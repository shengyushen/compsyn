// Benchmark "Huffman_random_9" written by ABC on Fri Nov 21 18:18:52 2014

module Huffman_random_9 ( clock, 
    in_0 , in_1 , in_2 , in_3 , in_4 , in_5 , in_6 , in_7 ,
    in_8 ,
    carestate, out  );
  input  clock;
  input  in_0 , in_1 , in_2 , in_3 , in_4 , in_5 , in_6 ,
    in_7 , in_8 ;
  output carestate, out;
  reg reg_0 , reg_1 , reg_2 , reg_3 , reg_4 , reg_5 , reg_6 ,
    reg_7 , reg_8 , counter_0 , counter_1 , counter_2 ,
    counter_3 , counter_4 ;
  wire n54_1, n64_1, n65, n66, n67, n68, n69_1, n70, n71, n72, n73, n74_1,
    n75, n76, n77, n78, n84_1, n85, n86, n87, n88, n89_1, n90, n91, n92,
    n93, n94, n96, n97, n24, n29, n34, n39, n44, n49, n54, n59, n64, n69,
    n74, n79, n84, n89;
  assign n54_1 = ~counter_0  & ~counter_1  & ~counter_2  & ~counter_3  & ~counter_4 ;
  assign n24 = n54_1 ? in_0  : reg_0 ;
  assign n29 = n54_1 ? in_1  : reg_1 ;
  assign n34 = n54_1 ? in_2  : reg_2 ;
  assign n39 = n54_1 ? in_3  : reg_3 ;
  assign n44 = n54_1 ? in_4  : reg_4 ;
  assign n49 = n54_1 ? in_5  : reg_5 ;
  assign n54 = n54_1 ? in_6  : reg_6 ;
  assign n59 = n54_1 ? in_7  : reg_7 ;
  assign n64 = n54_1 ? in_8  : reg_8 ;
  assign n64_1 = (~in_3  & ((~in_1  & in_5  & ((in_0  & ~in_2  & in_4  & (in_6  ^ in_7 )) | (~in_0  & in_2  & ~in_4  & in_6  & in_7 ))) | (~in_0  & in_1  & ~in_2  & ~in_6  & in_7  & in_4  & ~in_5 ))) | (~in_6  & in_7  & in_4  & ~in_5  & ~in_0  & in_1  & in_2  & in_3 ) | (in_4  & ((~in_0  & in_1  & in_2  & in_3  & ~in_5  & ~in_7  & (in_6  ^ in_8 )) | (in_0  & ~in_1  & ~in_2  & ~in_3  & in_5  & in_6  & in_7  & ~in_8 )));
  assign n65 = (in_3  & ((((in_0  & ~in_4  & ~in_5  & in_6 ) | (~in_0  & in_4  & in_5  & ~in_6 )) & (in_1  | (~in_1  & in_2 ))) | (~in_2  & ((in_0  & in_5  & (in_1  ^ in_4 )) | (~in_0  & ~in_1  & ~in_5 ) | (~in_4  & ((~in_0  & in_1  & in_5  & in_6 ) | (in_0  & ~in_1  & ~in_5  & ~in_6 ))))) | (~in_1  & in_2  & (((~in_4  ^ in_5 ) & (in_0  ^ in_6 )) | (~in_0  & in_4  & ~in_5  & ~in_6 ))))) | (~in_3  & (((in_1  ? (~in_4  ^ in_5 ) : (~in_4  & in_5 )) & (in_0  ? (in_2  ^ in_6 ) : (~in_2  & in_6 ))) | ((~in_4  ^ in_6 ) & ((~in_1  & ((~in_5  & (in_0  | (~in_0  & in_2 ))) | (~in_0  & ~in_2  & in_5 ))) | (~in_0  & in_1  & ~in_2  & ~in_5 ))) | (in_2  & ((in_5  & ((in_0  & in_6  & (~in_1  ^ in_4 )) | (~in_0  & in_1  & ~in_4  & ~in_6 ))) | (~in_0  & ~in_5  & (in_1  ? (in_4  & ~in_6 ) : (in_4  ^ in_6 ))))) | (~in_0  & ~in_2  & ((in_5  & in_6  & in_1  & ~in_4 ) | (~in_1  & in_4  & ~in_5  & ~in_6 ))))) | (~in_2  & (in_1  ? (in_4  ? (((~in_5  ^ in_7 ) & (in_0  ? (in_3  & in_6 ) : (~in_3  & ~in_6 ))) | (~in_5  & ((~in_6  & (in_0  ? ~in_7  : (in_3  & in_7 ))) | (in_6  & in_7  & ~in_0  & in_3 ))) | (~in_0  & in_3  & in_5  & in_6  & ~in_7 )) : ((in_7  & ((~in_0  & (in_3  ? ~in_5  : (in_5  & ~in_6 ))) | (in_5  & in_6  & in_0  & ~in_3 ))) | (in_0  & ~in_6  & ~in_7  & (~in_3  ^ ~in_5 )))) : (in_4  ? (((in_0  ^ in_5 ) & (in_3  ? (in_6  & ~in_7 ) : (~in_6  & in_7 ))) | (~in_3  & ~in_7  & (in_0  ? (in_5  & ~in_6 ) : (~in_5  & in_6 )))) : (((in_6  ^ in_7 ) & (in_0  ? (in_3  & in_5 ) : (~in_3  & ~in_5 ))) | (~in_0  & in_3  & in_5  & (~in_6  ^ in_7 )) | (in_0  & ~in_3  & ~in_5  & in_6  & in_7 ))))) | (in_2  & (in_0  ? ((~in_1  & in_3  & (in_4  ? (~in_5  & ~in_7 ) : (in_5  & in_7 ))) | (in_1  & ~in_3  & in_4  & ~in_5  & ~in_7 ) | (in_5  & (in_1  ? (~in_4  & (in_3  ? (~in_6  & ~in_7 ) : (~in_6  ^ in_7 ))) : (in_4  & (in_3  ? (in_6  & ~in_7 ) : (~in_6  & in_7 ))))) | (~in_1  & ~in_3  & in_4  & ~in_5  & ~in_6  & in_7 )) : (in_6  ? (((in_3  ? (in_4  & ~in_5 ) : (~in_4  & in_5 )) & (~in_1  ^ in_7 )) | (~in_7  & ((in_5  & ((~in_3  & in_4 ) | (in_3  & ~in_4 ) | (in_1  & in_3  & in_4 ))) | (~in_4  & ~in_5  & in_1  & ~in_3 )))) : ((~in_1  & ~in_4  & (in_3  ? (in_5  ^ in_7 ) : (in_5  & in_7 ))) | (in_1  & ~in_3  & in_4  & in_5  & in_7 ))))) | (~in_1  & (in_6  ? (in_0  ? ((~in_3  & ((in_4  & in_5  & (in_2  ? (~in_7  ^ ~in_8 ) : (in_7  & in_8 ))) | (~in_2  & ~in_4  & ~in_5  & ~in_7  & ~in_8 ))) | (~in_2  & in_3  & in_7  & (in_4  ? (~in_5  & ~in_8 ) : (in_5  ^ in_8 )))) : ((in_7  & ((in_3  & ((in_2  & ~in_8  & (~in_4  ^ ~in_5 )) | (~in_2  & in_4  & in_5  & in_8 ))) | (~in_2  & ~in_3  & ~in_5  & in_8 ))) | (~in_2  & in_3  & ~in_4  & in_5  & ~in_7  & in_8 ))) : (in_2  ? (((~in_3  ^ in_7 ) & ((in_0  & in_4  & ~in_5  & in_8 ) | (~in_0  & ~in_4  & in_5  & ~in_8 ))) | (in_5  & ((~in_7  & ((in_0  & (in_3  ? (~in_4  & ~in_8 ) : (in_4  & in_8 ))) | (~in_0  & ~in_3  & in_4  & ~in_8 ))) | (~in_0  & ~in_3  & in_4  & in_7  & in_8 )))) : ((in_8  & ((~in_0  & ((in_5  & in_7  & in_3  & in_4 ) | (~in_5  & ~in_7  & ~in_3  & ~in_4 ))) | (in_0  & in_3  & in_4  & ~in_5  & in_7 ))) | (in_5  & ~in_7  & ~in_8  & (~in_0  ^ ~in_4 )))))) | (in_1  & (in_0  ? (in_3  ? ((~in_6  & ((in_7  & ((~in_4  & (in_2  ? (in_5  ^ in_8 ) : (~in_5  & in_8 ))) | (in_5  & ~in_8  & ~in_2  & in_4 ))) | (~in_2  & in_4  & in_5  & ~in_7  & in_8 ))) | (~in_2  & in_4  & ~in_5  & in_6  & in_7  & ~in_8 )) : (in_2  ? ((~in_5  & ((in_4  & in_7  & (~in_6  ^ in_8 )) | (~in_4  & in_6  & ~in_7  & ~in_8 ))) | (~in_4  & in_5  & in_6  & ~in_7  & in_8 )) : (in_4  & ((~in_5  & in_7  & (~in_6  ^ in_8 )) | (in_5  & ~in_6  & ~in_7  & ~in_8 ))))) : (in_5  ? ((~in_8  & ((in_4  & ((in_6  & in_7  & (in_2  | (~in_2  & in_3 ))) | (~in_2  & ~in_3  & ~in_6  & ~in_7 ))) | (in_3  & ~in_4  & ~in_6  & ~in_7 ))) | (in_3  & ~in_4  & ~in_6  & in_7  & in_8 )) : ((in_8  & ((in_6  & ((in_3  & (in_2  ? (in_4  ^ in_7 ) : ~in_7 )) | (~in_4  & in_7  & in_2  & ~in_3 ))) | (in_2  & ~in_3  & ~in_4  & ~in_6  & in_7 ))) | (~in_2  & in_3  & ~in_4  & ~in_6  & ~in_7  & ~in_8 )))));
  assign n66 = ((in_3  ? (~in_4  & in_8 ) : (in_4  & ~in_8 )) & ((((~in_0  & (in_1  ? (~in_5  & ~in_7 ) : (in_5  & in_7 ))) | (in_0  & in_1  & in_5  & in_7 )) & (~in_2  ^ in_6 )) | (~in_5  & ((in_0  & in_1  & ~in_2  & in_6 ) | (~in_0  & ~in_1  & in_2  & ~in_6 ) | (in_0  & ~in_1  & ~in_2  & ~in_7 ) | (~in_0  & in_1  & in_2  & ~in_6  & in_7 ))) | (in_2  & in_5  & ((~in_6  & (in_0  ? (~in_1  ^ in_7 ) : (in_1  ^ in_7 ))) | (in_0  & in_6  & ~in_7 ))))) | (~in_5  & (in_1  ? (in_8  ? ((~in_6  & ((in_0  & (in_2  ? (in_3  & ~in_7 ) : (~in_3  & in_7 ))) | (~in_0  & in_2  & ~in_3  & ~in_7 ))) | (in_0  & ~in_2  & ~in_3  & in_6  & ~in_7 )) : ((in_3  & (in_2  ? ((~in_6  & (in_0  | (~in_0  & ~in_7 ))) | (~in_0  & in_6  & in_7 )) : (in_0  ? (~in_6  & in_7 ) : (in_6  & ~in_7 )))) | (in_2  & ~in_3  & in_6  & in_7 ))) : ((~in_8  & ((in_7  & ((in_3  & (in_0  ? (~in_2  ^ in_6 ) : (in_2  & ~in_6 ))) | (~in_0  & ~in_2  & ~in_3  & in_6 ))) | (in_0  & ~in_6  & ~in_7  & (in_2  ^ in_3 )))) | (in_6  & ~in_7  & in_8  & in_0  & ~in_2  & ~in_3 )))) | (in_5  & ((in_8  & (in_0  ? ((in_1  & ~in_3  & (in_2  ? (in_6  ^ in_7 ) : (~in_6  & in_7 ))) | (~in_1  & ~in_2  & in_3  & in_6  & in_7 )) : (in_2  ? ((in_6  & in_7  & in_1  & in_3 ) | (~in_6  & ~in_7  & ~in_1  & ~in_3 )) : ((~in_6  & (in_1  ? ~in_7  : (~in_3  & in_7 ))) | (in_6  & ~in_7  & ~in_1  & ~in_3 ))))) | (~in_2  & ~in_8  & ((in_3  & ~in_6  & (in_0  ? (in_1  & ~in_7 ) : in_7 )) | (~in_0  & ~in_1  & ~in_3  & in_6  & ~in_7 ))))) | (~in_2  & (in_7  ? ((~in_0  & in_4  & in_6  & (in_1  ? (~in_3  & in_5 ) : (~in_3  ^ ~in_5 ))) | (in_0  & ~in_1  & ~in_3  & ~in_4  & in_5  & ~in_6 )) : (in_0  ? (in_1  & ((~in_3  & ~in_4  & (~in_5  ^ in_6 )) | (in_5  & in_6  & in_3  & in_4 ))) : ((in_4  & ((in_1  & ~in_5  & (in_3  ^ in_6 )) | (in_5  & ~in_6  & ~in_1  & in_3 ))) | (~in_1  & in_3  & ~in_4  & ~in_5  & ~in_6 ))))) | (in_2  & ((~in_1  & ((~in_4  & ((~in_3  & ((~in_5  & (in_0  ? in_6  : (~in_6  & in_7 ))) | (in_6  & ~in_7  & ~in_0  & in_5 ))) | (in_0  & in_3  & ~in_5  & in_6  & ~in_7 ))) | (in_0  & in_3  & in_4  & in_5  & in_6  & in_7 ))) | (~in_0  & in_1  & ~in_3  & in_6  & ~in_7  & ~in_4  & in_5 ))) | (in_2  & (in_6  ? (in_7  ? (in_1  ? (in_3  ? ((~in_0  & (in_4  ? (~in_5  & in_8 ) : (in_5  & ~in_8 ))) | (in_0  & ~in_4  & in_5  & ~in_8 )) : (in_0  ? (~in_4  & (in_5  ^ in_8 )) : (in_4  & in_8 ))) : (in_4  & in_8  & (~in_3  ^ ~in_5 ))) : ((in_1  & ((in_0  & ~in_4  & in_5  & ~in_8 ) | (~in_0  & in_4  & ~in_5  & in_8 ) | (~in_4  & ~in_5  & (in_0  ? (~in_3  & in_8 ) : (in_3  & ~in_8 ))))) | (~in_4  & in_5  & ~in_8  & in_0  & ~in_1  & in_3 ))) : (in_1  ? (in_3  ? ((in_4  & ((in_0  & ~in_5  & in_7  & in_8 ) | (~in_0  & in_5  & ~in_7  & ~in_8 ))) | (~in_0  & ~in_4  & (in_5  ? (in_7  & ~in_8 ) : (~in_7  ^ ~in_8 )))) : (in_0  ? ((in_4  & in_8  & (in_5  ^ in_7 )) | (in_7  & ~in_8  & ~in_4  & in_5 )) : ((~in_4  & ~in_5  & ~in_8 ) | (in_4  & in_5  & ~in_7  & in_8 )))) : (~in_5  & (in_0  ? ((in_7  & (in_3  ? (~in_4  ^ ~in_8 ) : (~in_4  & ~in_8 ))) | (~in_3  & ~in_4  & ~in_7  & in_8 )) : ((in_3  & (in_4  ? in_8  : (~in_7  & ~in_8 ))) | (~in_3  & in_4  & ~in_7  & in_8 ))))))) | (~in_2  & (in_6  ? ((in_7  & ((in_4  & (in_0  ? ((~in_1  & (in_3  ? (in_5  ^ in_8 ) : (in_5  ^ ~in_8 ))) | (~in_5  & in_8  & in_1  & in_3 )) : (in_3  & (in_1  ? in_8  : (in_5  & ~in_8 ))))) | (in_0  & in_3  & ~in_4  & ~in_5  & ~in_8 ))) | (~in_4  & ~in_7  & ~in_8  & ((in_0  & ~in_5  & (~in_1  ^ ~in_3 )) | (~in_0  & ~in_1  & in_3  & in_5 )))) : (in_3  ? (in_1  ? ((in_5  & ((in_4  & (in_0  ? (in_7  & in_8 ) : (~in_7  ^ in_8 ))) | (in_0  & ~in_4  & (~in_7  ^ ~in_8 )))) | (in_0  & in_4  & ~in_5  & in_7  & in_8 )) : ((~in_4  & ((in_0  & in_8  & (in_5  ^ in_7 )) | (in_7  & ~in_8  & ~in_0  & ~in_5 ))) | (in_0  & in_4  & ~in_5  & ~in_7  & in_8 ))) : (in_0  ? (in_1  ? ((in_4  & in_5  & ~in_7  & in_8 ) | (~in_4  & in_7  & ~in_8 )) : (in_8  & (in_4  ? ~in_5  : (in_5  & ~in_7 )))) : (~in_7  & (in_1  ? (in_4  ? (~in_5  & in_8 ) : (in_5  & ~in_8 )) : (in_4  ? (in_5  & in_8 ) : (~in_5  & ~in_8 ))))))));
  assign n67 = (~in_3  & (in_1  ? (((in_0  ? (~in_2  & in_7 ) : (in_2  & ~in_7 )) & (in_5  | (~in_4  & ~in_5  & ~in_6 ))) | (in_6  & (in_0  ? ((~in_7  & (in_2  ? (~in_4  ^ in_5 ) : (~in_4  ^ ~in_5 ))) | (~in_4  & ~in_5  & in_7 )) : (in_4  & (in_2  ? (~in_5  | (in_5  & in_7 )) : (~in_5  & in_7 ))))) | (~in_4  & ~in_6  & ((in_0  & in_2  & in_7 ) | (~in_0  & ~in_2  & ~in_7 ) | (in_0  & ~in_5  & ~in_7 ) | (~in_0  & in_2  & in_5  & in_7 )))) : (((in_4  ^ in_7 ) & ((~in_2  & (in_0  ? ~in_6  : (in_5  & in_6 ))) | (~in_5  & in_6  & in_0  & in_2 ))) | (((~in_6  & in_7  & ~in_0  & in_4 ) | (in_6  & ~in_7  & in_0  & ~in_4 )) & (in_2  ^ in_5 )) | (in_2  & ((in_6  & ((~in_0  & (in_4  ? (~in_5  ^ in_7 ) : (~in_5  & ~in_7 ))) | (in_0  & ~in_4  & in_5  & ~in_7 ))) | (~in_5  & ~in_6  & (~in_7  | (in_0  & in_4  & in_7 )))))))) | (in_3  & ((~in_7  & (((~in_1  ^ in_4 ) & (in_2  ? (~in_5  & ~in_6 ) : (in_5  & in_6 ))) | (~in_4  & ~in_5  & ~in_6  & in_1  & in_2 ))) | (in_5  & in_6  & in_7  & in_1  & in_2  & ~in_4 ) | (~in_1  & in_7  & ((in_0  & in_2  & in_6 ) | (~in_4  & ~in_6  & ~in_0  & ~in_2 ))) | (~in_0  & in_1  & ~in_2  & ~in_7  & (in_4  ^ in_6 )) | (~in_1  & (in_0  ? ((~in_7  & (in_4  ^ in_6 ) & (in_2  ^ ~in_5 )) | (in_5  & in_7  & (in_2  ? (in_4  & ~in_6 ) : (~in_4  & in_6 )))) : ((in_6  & ((~in_7  & (in_2  ? (~in_4  ^ in_5 ) : (in_4  & ~in_5 ))) | (~in_5  & in_7  & ~in_2  & ~in_4 ))) | (~in_4  & ~in_6  & (in_2  ? (in_5  & in_7 ) : (~in_5  & ~in_7 )))))) | (in_1  & (in_4  ? (~in_6  & in_7  & (in_0  ? ~in_5  : (in_2  & in_5 ))) : (in_6  ? ((in_5  & in_7  & in_0  & ~in_2 ) | (~in_0  & in_2  & ~in_5  & ~in_7 )) : (((in_2  ^ ~in_7 ) & (in_0  ^ ~in_5 )) | (in_5  & ~in_7  & in_0  & in_2 ))))))) | (~in_0  & (in_1  ? (in_3  & ((in_7  & ((in_6  & (in_4  ? (in_5  ^ ~in_8 ) : (~in_5  & ~in_8 ))) | (~in_4  & in_5  & ~in_6  & ~in_8 ))) | (~in_4  & in_5  & ~in_6  & ~in_7  & in_8 ))) : (~in_3  & ((in_4  & in_5  & ~in_6  & ~in_7  & in_8 ) | (~in_4  & ~in_5  & in_6  & in_7  & ~in_8 ))))) | (in_0  & (in_5  ? ((~in_1  & in_8  & ((in_6  & in_7  & ~in_3  & in_4 ) | (~in_6  & ~in_7  & in_3  & ~in_4 ))) | (in_1  & in_3  & ~in_4  & in_6  & ~in_7  & ~in_8 )) : (~in_6  & ((in_7  & ((in_1  & (in_3  ? (~in_4  & ~in_8 ) : (in_4  & in_8 ))) | (in_4  & ~in_8  & ~in_1  & in_3 ))) | (in_1  & ~in_3  & in_4  & ~in_7  & ~in_8 ))))) | (((~in_6  & ((~in_5  & ((in_2  & in_7  & (in_3  ^ in_8 )) | (~in_2  & ~in_3  & ~in_7  & in_8 ))) | (~in_2  & ~in_3  & in_5  & ~in_7  & in_8 ))) | (in_6  & ~in_7  & in_8  & in_2  & in_3  & ~in_5 )) & (in_0  ? (~in_1  & ~in_4 ) : (in_1  & in_4 ))) | (~in_1  & (in_2  ? (in_7  ? ((~in_0  & ((in_5  & ((in_8  & (in_3  ? (in_4  ^ in_6 ) : (~in_4  & ~in_6 ))) | (~in_3  & in_4  & ~in_6  & ~in_8 ))) | (in_3  & ~in_5  & in_6  & (~in_4  ^ in_8 )))) | (in_0  & ~in_3  & in_4  & ~in_5  & in_6  & ~in_8 )) : ((~in_0  & ((~in_3  & ~in_4  & in_5  & in_8 ) | (in_3  & in_4  & ~in_5  & ~in_8 ))) | (in_0  & ~in_3  & in_4  & in_5  & ~in_8 ) | (~in_0  & in_3  & ~in_4  & in_5  & ~in_6  & in_8 ))) : (((~in_4  ^ in_7 ) & ((in_0  & ~in_3  & ~in_5  & in_6  & in_8 ) | (~in_0  & in_3  & in_5  & ~in_6  & ~in_8 ))) | (in_3  & (in_4  ? ((in_8  & (((in_5  ^ in_7 ) & (~in_0  ^ in_6 )) | (in_6  & in_7  & in_0  & in_5 ))) | (~in_0  & in_5  & in_6  & in_7  & ~in_8 )) : (in_6  & ~in_8  & (in_0  ? (~in_5  & in_7 ) : (~in_5  ^ in_7 ))))) | (~in_0  & ~in_3  & ~in_8  & ((~in_6  & (in_4  ? (~in_5  & ~in_7 ) : (~in_5  ^ in_7 ))) | (in_4  & in_6  & in_7 )))))) | (in_1  & (in_5  ? (in_4  ? ((~in_6  & ((in_3  & ((~in_2  & (in_0  ? (~in_7  ^ in_8 ) : (in_7  & ~in_8 ))) | (~in_0  & in_2  & ~in_7  & in_8 ))) | (in_0  & ~in_3  & ~in_7  & (in_2  ^ in_8 )))) | (~in_2  & in_6  & in_8  & (in_0  ? (in_3  & in_7 ) : (~in_3  & ~in_7 )))) : ((in_6  & ((~in_3  & ((in_0  & in_2  & (~in_7  ^ in_8 )) | (in_7  & in_8  & ~in_0  & ~in_2 ))) | (~in_0  & ~in_2  & in_3  & in_7  & ~in_8 ))) | (in_0  & ~in_2  & in_3  & ~in_6  & in_7  & ~in_8 ))) : ((~in_8  & ((in_4  & ((~in_2  & (in_0  ? (in_3  ? (~in_6  & ~in_7 ) : (in_6  & in_7 )) : (in_6  & ~in_7 ))) | (~in_0  & in_2  & ~in_3  & ~in_6  & ~in_7 ))) | (~in_0  & in_2  & ~in_3  & ~in_4  & in_7 ))) | (in_0  & ~in_2  & in_3  & in_4  & in_6  & in_7  & in_8 ))));
  assign n68 = ((in_1  ^ in_4 ) & (((in_3  ? (in_5  & ~in_6 ) : (~in_5  & in_6 )) & ((~in_0  & in_7  & ~in_8 ) | (~in_7  & in_8  & in_0  & in_2 ))) | (in_0  & (in_3  ? ((in_5  & ((~in_2  & ~in_7  & in_8 ) | (in_2  & in_7  & ~in_8 ) | (in_6  & in_7  & in_8 ))) | (in_2  & ~in_5  & (in_6  ? (~in_7  ^ in_8 ) : (~in_7  & ~in_8 )))) : ((~in_5  & (in_2  ? (~in_6  & (~in_7  | (in_7  & ~in_8 ))) : (in_6  ? (in_7  & ~in_8 ) : (~in_7  & in_8 )))) | (in_2  & in_5  & (in_6  ? (~in_7  ^ in_8 ) : in_7 ))))) | (~in_0  & (in_2  ? ((in_3  & ((~in_7  & ((~in_6  & in_8 ) | (in_6  & ~in_8 ) | (in_5  & in_6  & in_8 ))) | (in_5  & in_6  & in_7  & in_8 ))) | (~in_3  & in_5  & in_6  & in_7  & in_8 )) : (in_8  & ((~in_3  & (in_5  ? (~in_6  ^ in_7 ) : (in_6  & ~in_7 ))) | (in_6  & in_7  & in_3  & ~in_5 ))))))) | (in_8  & ((((~in_6  & in_7  & ~in_3  & in_4 ) | (in_6  & ~in_7  & in_3  & ~in_4 )) & ((in_5  & (in_0  ? (in_1  & in_2 ) : (~in_1  ^ ~in_2 ))) | (in_0  & ~in_5  & (in_1  ^ ~in_2 )))) | (~in_1  & ~in_4  & ((~in_5  & ((~in_0  & (in_2  ? (~in_3  & ~in_7 ) : in_3 )) | (~in_3  & in_7  & in_0  & ~in_2 ))) | (in_3  & in_5  & ((in_0  & ~in_2  & in_7 ) | (in_0  & ~in_7 ) | (~in_0  & in_7 ))))) | (in_1  & in_4  & ((~in_0  & in_2  & in_3  & in_7 ) | (~in_3  & ~in_7  & in_0  & ~in_2 ) | (~in_0  & ((in_5  & (in_2  ? (in_3  ^ in_7 ) : (in_3  & ~in_7 ))) | (~in_2  & ~in_3  & ~in_5  & ~in_7 ))) | (in_0  & ~in_2  & in_3  & ~in_5  & in_7 ))) | (in_4  & (in_2  ? (in_5  ? ((in_0  & ~in_1  & in_3  & ~in_6  & in_7 ) | (~in_0  & in_1  & ~in_3  & in_6  & ~in_7 )) : ((in_3  & (((in_0  ^ in_6 ) & (in_1  ^ in_7 )) | (~in_0  & ~in_1  & in_6  & ~in_7 ))) | (in_1  & ~in_3  & (in_0  ? (~in_6  ^ in_7 ) : (in_6  & in_7 ))))) : (in_5  ? (in_0  ? (in_6  & (in_1  ? in_3  : (~in_3  & ~in_7 ))) : (in_1  ? (in_3  ? (in_6  & in_7 ) : (~in_6  & ~in_7 )) : (in_3  ? (~in_6  & in_7 ) : (in_6  & ~in_7 )))) : (((in_0  ^ in_6 ) & (in_1  ? (~in_3  & in_7 ) : (in_3  & ~in_7 ))) | (in_6  & ((in_0  & ~in_1  & ~in_3 ) | (in_1  & in_3  & (~in_0  ^ ~in_7 )))) | (~in_0  & in_3  & ~in_6  & (in_1  ^ in_7 )))))) | (~in_4  & (in_5  ? (in_0  ? (~in_2  & ~in_3  & (in_1  ? (in_6  & in_7 ) : ~in_6 )) : ((~in_2  & ((in_3  & (in_1  ? (~in_6  ^ in_7 ) : (~in_6  & ~in_7 ))) | (~in_6  & in_7  & ~in_1  & ~in_3 ))) | (~in_1  & in_2  & ~in_3  & (in_6  ^ in_7 )))) : (((in_2  ^ ~in_7 ) & ((in_0  & ~in_1  & ~in_3  & in_6 ) | (~in_0  & in_1  & in_3  & ~in_6 ))) | (~in_0  & ((~in_3  & ((in_1  & (in_2  ? (in_6  & ~in_7 ) : (~in_6  & in_7 ))) | (~in_6  & ~in_7  & ~in_1  & ~in_2 ))) | (~in_1  & in_2  & in_3  & in_6 ))) | (in_0  & in_6  & in_7  & (in_1  ? (in_2  ^ in_3 ) : (in_2  & in_3 )))))))) | (~in_8  & (((in_3  ^ in_6 ) & (in_0  ? (in_4  & ((~in_5  & ((~in_1  & ~in_2  & ~in_7 ) | (in_7  & (in_1  | (~in_1  & in_2 ))))) | (in_5  & ~in_7  & ~in_1  & ~in_2 ))) : (in_7  ? ((in_4  & in_5  & in_1  & in_2 ) | (~in_4  & ~in_5  & ~in_1  & ~in_2 )) : ((in_5  & (in_1  ? (~in_2  & in_4 ) : (in_2  ^ ~in_4 ))) | (in_1  & in_2  & ~in_5 ))))) | ((in_5  ? (in_6  & in_7 ) : (~in_6  & ~in_7 )) & ((~in_2  & ((~in_4  & (in_0  ? ~in_1  : (in_1  & in_3 ))) | (~in_0  & in_1  & in_3  & in_4 ))) | (in_0  & ~in_1  & in_2  & ~in_3  & ~in_4 ))) | (~in_0  & (in_4  ? (~in_7  & (in_1  ? (in_2  ? (~in_3  & ~in_6 ) : (in_3  & in_6 )) : (~in_2  & in_6 ))) : ((in_2  & in_3  & (in_1  ? (in_6  & in_7 ) : ~in_7 )) | (~in_3  & ~in_6  & in_7  & ~in_1  & ~in_2 )))) | (in_0  & ((in_1  & ~in_2  & ((~in_7  & (in_3  ? in_4  : (~in_4  & ~in_6 ))) | (~in_6  & in_7  & ~in_3  & ~in_4 ))) | (~in_1  & in_2  & in_3  & ~in_4  & in_6  & ~in_7 ))) | (~in_1  & (in_0  ? ((~in_2  & ~in_3  & ~in_4  & ~in_5  & in_7 ) | (in_2  & in_3  & in_4  & in_5  & ~in_7 ) | (in_3  & in_6  & ((~in_2  & (in_4  ? in_5  : (~in_5  & in_7 ))) | (~in_5  & in_7  & in_2  & in_4 )))) : (in_4  ? (in_7  & (in_2  ? (in_3  ? (~in_5  & ~in_6 ) : (in_5  & in_6 )) : (in_3  & ~in_5 ))) : (in_2  ? (in_7  & (in_3  ? (~in_5  & in_6 ) : (in_5  ^ in_6 ))) : (~in_7  & (in_3  ? (in_5  & in_6 ) : (~in_5  & ~in_6 ))))))) | (in_1  & ((~in_2  & (in_0  ? ((in_3  & ~in_4  & (in_5  ? (~in_6  & in_7 ) : (in_6  & ~in_7 ))) | (~in_3  & in_4  & ~in_5  & ~in_6  & ~in_7 )) : ((~in_3  & ((in_4  & (in_5  ? ~in_6  : (in_6  & in_7 ))) | (~in_6  & in_7  & ~in_4  & ~in_5 ))) | (~in_5  & in_6  & in_7  & in_3  & in_4 )))) | (~in_0  & in_2  & ((in_3  & in_4  & in_5  & in_6 ) | (~in_5  & ~in_6  & in_7  & ~in_3  & ~in_4 )))))));
  assign n69_1 = 1'b0;
  assign n70 = counter_4  | n69_1;
  assign n71 = counter_3  | n70;
  assign n72 = counter_2  | n71;
  assign n73 = counter_1  | n72;
  assign n74_1 = counter_0  ^ ~n73;
  assign n75 = counter_1  ^ ~n72;
  assign n76 = counter_2  ^ ~n71;
  assign n77 = counter_3  ^ ~n70;
  assign n78 = counter_4  ^ ~n69_1;
  assign n69 = n54_1 ? n64_1 : n74_1;
  assign n74 = n54_1 ? n65 : n75;
  assign n79 = n54_1 ? n66 : n76;
  assign n84 = n54_1 ? n67 : n77;
  assign n89 = n54_1 ? n68 : n78;
  assign n84_1 = in_0  ^ ~reg_0 ;
  assign n85 = in_1  ^ ~reg_1 ;
  assign n86 = in_2  ^ ~reg_2 ;
  assign n87 = in_3  ^ ~reg_3 ;
  assign n88 = in_4  ^ ~reg_4 ;
  assign n89_1 = in_5  ^ ~reg_5 ;
  assign n90 = in_6  ^ ~reg_6 ;
  assign n91 = in_7  ^ ~reg_7 ;
  assign n92 = in_8  ^ ~reg_8 ;
  assign n93 = n92 & n91 & n90 & n89_1 & n88 & n87 & n86 & n84_1 & n85;
  assign n94 = in_0  & in_1  & in_2  & in_3  & in_4  & (in_5  | (~in_5  & in_6 ));
  assign carestate = n54_1 ? ~n94 : n93;
  assign n96 = in_0  & (in_1  | (~in_1  & in_2 ) | (in_3  & in_4  & ~in_1  & ~in_2 ) | (~in_1  & ~in_2  & in_3  & ~in_4  & in_5 ) | (~in_1  & ~in_2  & in_3  & in_6  & in_7  & ~in_4  & ~in_5 ) | (in_3  & ~in_4  & ~in_1  & ~in_2  & ~in_5  & in_6  & ~in_7  & in_8 ));
  assign n97 = ((reg_7  ^ reg_8 ) & ((~counter_1  & (counter_3  ? ((~counter_0  & ((((~reg_0  & ~reg_2  & ~reg_4  & reg_6 ) | (reg_0  & reg_2  & reg_4  & ~reg_6 )) & ((reg_1  & ((counter_2  & reg_3  & ~reg_5 ) | (~counter_2  & counter_4  & ~reg_3  & reg_5 ))) | (counter_2  & ~counter_4  & ~reg_1  & ~reg_3  & reg_5 ))) | (counter_2  & (counter_4  ? (~reg_2  & ~reg_3  & ~reg_5  & (reg_0  ? reg_4  : (reg_1  & ~reg_4 ))) : ((~reg_3  & ((~reg_0  & reg_1  & ~reg_4  & reg_5 ) | (reg_0  & ~reg_1  & reg_4  & ~reg_5 ) | (~reg_0  & reg_2  & reg_4  & (~reg_1  ^ reg_5 )))) | (~reg_0  & reg_1  & reg_2  & reg_3  & ~reg_4 )))) | (~counter_2  & ((~reg_3  & ((~reg_0  & reg_2  & ((counter_4  & reg_1  & (~reg_4  ^ reg_5 )) | (~counter_4  & ~reg_1  & ~reg_4  & ~reg_5 ))) | (~counter_4  & reg_0  & reg_1  & ~reg_2  & reg_4  & reg_5 ))) | (counter_4  & ~reg_1  & ~reg_2  & reg_3  & ~reg_5  & (~reg_0  ^ reg_4 )))) | ((~reg_2  ^ ~reg_6 ) & ((reg_1  & ((~reg_4  & reg_5  & ((counter_2  & (counter_4  ? (~reg_0  & ~reg_3 ) : (reg_0  & reg_3 ))) | (~reg_0  & reg_3  & ~counter_2  & ~counter_4 ))) | (~counter_2  & ~counter_4  & ~reg_0  & ~reg_3  & reg_4  & ~reg_5 ))) | (counter_2  & counter_4  & reg_0  & ~reg_1  & (reg_3  ? (reg_4  & reg_5 ) : (~reg_4  & ~reg_5 ))))) | ((reg_1  ^ reg_2 ) & ((~reg_0  & reg_6  & ((~counter_2  & ((~counter_4  & reg_3  & reg_4  & reg_5 ) | (counter_4  & ~reg_3  & ~reg_4  & ~reg_5 ))) | (counter_2  & counter_4  & ~reg_3  & reg_4  & ~reg_5 ))) | (counter_2  & ~counter_4  & reg_0  & ~reg_3  & ~reg_4  & ~reg_6 ))) | (~reg_1  & (((~reg_2  ^ reg_6 ) & ((reg_0  & ((counter_2  & ((counter_4  & ~reg_3  & reg_4  & reg_5 ) | (~counter_4  & reg_3  & ~reg_4  & ~reg_5 ))) | (~counter_2  & counter_4  & reg_3  & ~reg_4  & ~reg_5 ))) | (reg_3  & ~reg_4  & ~reg_5  & ~counter_2  & ~counter_4  & ~reg_0 ))) | ((~reg_4  ^ reg_6 ) & ((~reg_0  & reg_3  & reg_5  & (counter_2  ? (counter_4  & reg_2 ) : (~counter_4  ^ reg_2 ))) | (~counter_2  & ~counter_4  & reg_0  & ~reg_3  & ~reg_5 ))) | (reg_3  & (counter_4  ? (~reg_2  & ((~counter_2  & ((reg_5  & (reg_0  ? reg_6  : (~reg_4  & ~reg_6 ))) | (~reg_5  & reg_6  & ~reg_0  & reg_4 ))) | (counter_2  & reg_0  & ~reg_4  & reg_5  & reg_6 ))) : (reg_0  ? (reg_6  & (((reg_2  ^ reg_4 ) & (~counter_2  ^ reg_5 )) | (~counter_2  & (reg_2  ? (reg_4  & ~reg_5 ) : (~reg_4  & reg_5 ))))) : (~reg_6  & ((~counter_2  & (reg_2  ? (~reg_4  & reg_5 ) : (reg_4  & ~reg_5 ))) | (counter_2  & reg_2  & reg_4  & reg_5 )))))) | (~reg_3  & ((~reg_6  & ((~counter_4  & ((counter_2  & reg_0  & ~reg_2  & ~reg_4  & reg_5 ) | (~counter_2  & ~reg_0  & reg_2  & reg_4  & ~reg_5 ))) | (~counter_2  & counter_4  & ~reg_0  & ~reg_5  & (~reg_2  | (reg_2  & reg_4 ))))) | (counter_4  & reg_0  & reg_6  & ((counter_2  & ~reg_4  & reg_5 ) | (~counter_2  & reg_2  & reg_4  & ~reg_5 ))))))) | (reg_1  & (((counter_2  ? (~counter_4  & ~reg_5 ) : (counter_4  & reg_5 )) & ((~reg_0  & ~reg_2  & ~reg_3  & reg_4  & reg_6 ) | (reg_0  & reg_2  & reg_3  & ~reg_4  & ~reg_6 ))) | (reg_5  & (reg_2  ? (reg_4  ? (reg_6  & ((~reg_0  & (counter_2  ^ ~counter_4 )) | (reg_0  & ~reg_3  & ~counter_2  & ~counter_4 ))) : ((~reg_6  & ((counter_4  & (counter_2  ? reg_3  : (~reg_0  & ~reg_3 ))) | (~counter_2  & ~counter_4  & reg_0 ))) | (counter_2  & ~counter_4  & reg_0  & ~reg_3  & reg_6 ))) : (~reg_6  & (counter_4  ? (reg_0  & reg_3  & (~counter_2  | (counter_2  & ~reg_4 ))) : ((reg_4  & (counter_2  ? (reg_0  ^ ~reg_3 ) : (reg_0  & reg_3 ))) | (~counter_2  & reg_0  & reg_3  & ~reg_4 )))))) | (~reg_5  & (counter_2  ? (~counter_4  & ((~reg_0  & ((reg_2  & ~reg_3  & reg_4  & reg_6 ) | (~reg_2  & reg_3  & ~reg_4  & ~reg_6 ))) | (reg_0  & ~reg_2  & ~reg_3  & reg_4  & ~reg_6 ))) : ((reg_0  & ((reg_2  & ((reg_3  & (counter_4  ? ~reg_6  : (~reg_4  & reg_6 ))) | (~counter_4  & ~reg_3  & ~reg_4  & ~reg_6 ))) | (~counter_4  & ~reg_2  & reg_3  & reg_4  & ~reg_6 ))) | (~counter_4  & ~reg_0  & ~reg_4  & (reg_2  ? (~reg_3  & reg_6 ) : (reg_3  & ~reg_6 )))))))))) | (counter_0  & ~counter_2  & ~counter_4  & ~reg_0  & reg_1  & reg_2  & reg_3  & reg_4  & ~reg_5  & ~reg_6 )) : ((~counter_2  & ((((reg_0  & ~reg_1  & ~reg_2  & ~reg_3  & reg_5  & reg_6 ) | (~reg_0  & reg_1  & reg_2  & reg_3  & ~reg_5  & ~reg_6 )) & (counter_0  ? (~counter_4  & reg_4 ) : (counter_4  & ~reg_4 ))) | (counter_4  & ((reg_4  & ((~reg_0  & ((reg_3  & ((~counter_0  & ((reg_6  & (reg_2  ^ reg_5 )) | (reg_1  & ~reg_2  & reg_5  & ~reg_6 ))) | (counter_0  & reg_1  & reg_2  & ~reg_5  & ~reg_6 ))) | (~counter_0  & ~reg_1  & ~reg_3  & reg_6  & (reg_2  | (~reg_2  & reg_5 ))))) | (~counter_0  & reg_0  & (reg_2  ? ((reg_6  & (reg_1  ? ~reg_3  : (reg_3  & reg_5 ))) | (reg_1  & ~reg_3  & ~reg_5  & ~reg_6 )) : (reg_1  ? (~reg_5  & (~reg_3  ^ reg_6 )) : (reg_5  & (reg_3  ^ reg_6 ))))))) | (~counter_0  & ~reg_4  & (reg_5  ? ((~reg_0  & reg_2  & reg_3  & reg_6 ) | (reg_0  & ~reg_2  & ~reg_3  & ~reg_6 ) | (~reg_1  & ~reg_3  & (~reg_0  ^ reg_2 ) & reg_6 )) : ((~reg_3  & ((reg_0  & (reg_1  ? reg_6  : (reg_2  & ~reg_6 ))) | (~reg_0  & ~reg_1  & ~reg_2  & reg_6 ))) | (reg_0  & reg_1  & ~reg_2  & reg_3  & ~reg_6 )))))))) | (~counter_0  & counter_2  & (reg_2  ? (reg_1  ? (((reg_4  ^ reg_5 ) & (((reg_0  ^ ~reg_3 ) & ~reg_6 ) | (~counter_4  & ~reg_0  & ~reg_3  & reg_6 ))) | (~counter_4  & ~reg_3  & (reg_0  ? (~reg_4  ^ reg_5 ) : (reg_4  & reg_5 ))) | (counter_4  & reg_0  & reg_3  & ~reg_4  & ~reg_5 ) | (~reg_4  & ((reg_0  & ((reg_5  & (~reg_3  ^ reg_6 )) | (~counter_4  & reg_3  & ~reg_5  & reg_6 ))) | (~counter_4  & ~reg_0  & reg_3  & reg_5  & ~reg_6 )))) : (((counter_4  ? (~reg_0  & reg_5 ) : ~reg_5 ) & (reg_3  ? (reg_4  & ~reg_6 ) : (~reg_4  & reg_6 ))) | (counter_4  & reg_0  & ~reg_5  & (reg_3  ^ reg_4 )) | (~counter_4  & ~reg_0  & reg_3  & reg_4  & reg_5 ) | (reg_4  & (counter_4  ? ((~reg_0  & reg_3  & ~reg_5  & reg_6 ) | (reg_0  & ~reg_3  & reg_5  & ~reg_6 )) : ((reg_0  & reg_5  & (~reg_3  ^ reg_6 )) | (~reg_0  & ~reg_3  & ~reg_5  & ~reg_6 )))) | (~counter_4  & reg_0  & ~reg_3  & ~reg_4  & ~reg_5  & ~reg_6 ))) : ((~counter_4  & ~reg_0  & reg_6  & (reg_1  ? reg_5  : (reg_3  & ~reg_5 ))) | (counter_4  & reg_0  & reg_1  & ~reg_3  & ~reg_5  & ~reg_6 ) | (~reg_1  & (((~counter_4  ^ reg_0 ) & (reg_3  ? (reg_4  ? (reg_5  & reg_6 ) : (~reg_5  & ~reg_6 )) : (~reg_6  & (reg_4  ^ reg_5 )))) | (reg_4  & ((~reg_5  & ((reg_6  & (counter_4  ? reg_3  : (~reg_0  & ~reg_3 ))) | (~counter_4  & reg_0  & ~reg_3  & ~reg_6 ))) | (reg_0  & reg_3  & reg_5  & ~reg_6 ))) | (reg_0  & ~reg_4  & ((~counter_4  & reg_3  & (~reg_5  ^ reg_6 )) | (counter_4  & ~reg_3  & ~reg_5  & reg_6 ))))) | (reg_1  & ((reg_3  & ((~reg_5  & (counter_4  ? (~reg_4  & (~reg_0  | (reg_0  & reg_6 ))) : (reg_0  ? (reg_4  ^ reg_6 ) : (reg_4  & reg_6 )))) | (counter_4  & reg_5  & (reg_0  ? (~reg_4  ^ reg_6 ) : (~reg_4  & reg_6 ))))) | (counter_4  & ~reg_0  & ~reg_3  & reg_4  & ~reg_5  & ~reg_6 ))))))))) | (~counter_0  & counter_1  & (reg_0  ? (reg_2  ? (reg_3  ? ((~counter_2  & ((~reg_6  & ((~reg_4  & ((reg_1  & reg_5  & (counter_3  | (~counter_3  & ~counter_4 ))) | (~counter_3  & counter_4  & ~reg_1  & ~reg_5 ))) | (~counter_4  & ~reg_1  & reg_4  & reg_5 ))) | (~counter_3  & ~reg_4  & ~reg_5  & (counter_4  ^ reg_1 ) & reg_6 ))) | (counter_2  & ~counter_3  & counter_4  & ~reg_5  & reg_6  & ~reg_1  & ~reg_4 )) : ((reg_1  & ((reg_5  & (((reg_4  ^ reg_6 ) & (counter_2  ? (~counter_3  & ~counter_4 ) : (counter_3  & counter_4 ))) | (~counter_2  & counter_4  & reg_4  & (~counter_3  ^ reg_6 )))) | (~counter_2  & ~reg_5  & ~reg_6  & ((~reg_4  & (~counter_3  | (counter_3  & counter_4 ))) | (~counter_3  & ~counter_4  & reg_4 ))))) | (~counter_2  & ~counter_3  & ~reg_1  & ~reg_5  & (reg_4  | (~reg_4  & ~reg_6 ))))) : (reg_5  ? ((counter_3  & ((~counter_4  & ~reg_1  & ~reg_3  & reg_4  & reg_6 ) | (counter_4  & reg_1  & reg_3  & ~reg_4  & ~reg_6 ))) | (~counter_3  & ((counter_4  & ~reg_1  & ~reg_3  & reg_4  & reg_6 ) | (~counter_4  & reg_1  & reg_3  & ~reg_4  & ~reg_6 ))) | (~reg_1  & ((~reg_3  & ((reg_4  & ((counter_3  & (counter_2  ? (counter_4  & reg_6 ) : (~counter_4  & ~reg_6 ))) | (~counter_2  & ~counter_3  & (~counter_4  | (counter_4  & ~reg_6 ))))) | (~counter_2  & ~counter_3  & ~reg_4  & reg_6 ))) | (~counter_2  & ~counter_3  & ~counter_4  & reg_3  & reg_4  & reg_6 ))) | (~counter_2  & ~counter_3  & ~counter_4  & reg_1  & reg_3  & reg_4  & ~reg_6 )) : ((~reg_4  & (((~reg_1  ^ reg_6 ) & ((~counter_2  & (counter_3  ? (~counter_4  & ~reg_3 ) : reg_3 )) | (counter_2  & ~counter_3  & ~counter_4  & reg_3 ))) | (~counter_2  & ~reg_1  & ~reg_6  & (counter_3  ? reg_3  : (counter_4  & ~reg_3 ))))) | (~reg_1  & ~reg_3  & reg_4  & reg_6  & ((~counter_2  & counter_3 ) | (counter_2  & ~counter_3 ) | (~counter_2  & ~counter_3  & counter_4 )))))) : (reg_4  ? (reg_1  ? (counter_4  ? ((~counter_2  & ((reg_2  & reg_5  & (reg_3  ^ reg_6 )) | (~reg_2  & ~reg_3  & ~reg_5  & ~reg_6 ) | (~counter_3  & reg_6  & (reg_2  ? (reg_3  & reg_5 ) : ~reg_3 )))) | (counter_2  & ~counter_3  & reg_2  & reg_3  & ~reg_5  & reg_6 )) : (counter_3  ? ((~reg_5  & (counter_2  ? (reg_2  ? (reg_3  & reg_6 ) : (~reg_3  & ~reg_6 )) : (~reg_3  & ~reg_6 ))) | (~counter_2  & reg_3  & reg_5  & ~reg_6 )) : (reg_2  & ((~counter_2  & (reg_3  ? (reg_5  & reg_6 ) : (~reg_5  ^ reg_6 ))) | (counter_2  & ~reg_3  & ~reg_5  & ~reg_6 ))))) : ((reg_2  & ~reg_6  & ((~reg_5  & ((~counter_4  & (counter_2  ^ counter_3 )) | (~counter_2  & counter_4  & (counter_3  ^ reg_3 )))) | (~counter_2  & ~counter_3  & ~counter_4  & reg_3  & reg_5 ))) | (~counter_2  & ~counter_3  & counter_4  & ~reg_2  & ~reg_3  & reg_5  & reg_6 ))) : ((~counter_3  & ((~reg_1  & (counter_4  ? ((~counter_2  & ((~reg_6  & (reg_2  ? (~reg_3  ^ reg_5 ) : (reg_3  & ~reg_5 ))) | (reg_2  & ~reg_3  & ~reg_5  & reg_6 ))) | (counter_2  & reg_2  & ~reg_3  & reg_5  & reg_6 )) : (counter_2  ? ((reg_2  & ~reg_3  & reg_5  & reg_6 ) | (~reg_2  & reg_3  & ~reg_5  & ~reg_6 )) : (reg_6  & (reg_2  ? ~reg_5  : (reg_3  & reg_5 )))))) | (~counter_2  & reg_1  & ~reg_2  & ~reg_5  & reg_6  & (~counter_4  | (counter_4  & reg_3 ))))) | (~counter_2  & counter_3  & ((reg_1  & reg_5  & ((counter_4  & ~reg_2  & reg_3  & reg_6 ) | (~counter_4  & reg_2  & ~reg_3  & ~reg_6 ))) | (~counter_4  & ~reg_1  & reg_3  & ~reg_5  & (~reg_2  ^ reg_6 )))))))))) | (~counter_1  & ((~reg_3  & (((counter_4  ? (reg_6  & ~reg_7 ) : (~reg_6  & reg_7 )) & ((~counter_0  & reg_1  & ~reg_5  & ((~counter_2  & counter_3  & (~reg_0  ^ reg_2 ) & reg_4 ) | (counter_2  & ~counter_3  & ~reg_0  & reg_2  & ~reg_4 ))) | (~counter_3  & reg_0  & counter_0  & ~counter_2  & ~reg_1  & ~reg_2  & reg_4  & reg_5 ))) | (~counter_0  & (((reg_0  ^ reg_6 ) & ((~reg_2  & ((reg_7  & ((counter_2  & ~counter_4  & ((~counter_3  & (reg_1  ? (reg_4  & ~reg_5 ) : (~reg_4  & reg_5 ))) | (counter_3  & reg_1  & reg_4  & reg_5 ))) | (~counter_2  & ~counter_3  & counter_4  & reg_1  & ~reg_4  & ~reg_5 ))) | (~counter_2  & counter_3  & counter_4  & ~reg_1  & reg_4  & ~reg_7 ))) | (~counter_4  & ~reg_1  & counter_2  & ~counter_3  & reg_2  & ~reg_4  & reg_5  & ~reg_7 ))) | (counter_2  & (((reg_6  ^ reg_7 ) & ((counter_3  & ((counter_4  & reg_1  & reg_4  & (reg_0  ? (reg_2  & ~reg_5 ) : (~reg_2  & reg_5 ))) | (~counter_4  & reg_0  & ~reg_1  & ~reg_2  & ~reg_4  & ~reg_5 ))) | (~counter_3  & counter_4  & reg_0  & reg_1  & ~reg_2  & ~reg_4  & reg_5 ))) | (~reg_4  & (counter_4  ? (counter_3  ? (reg_0  ? ((reg_1  & (reg_2  ? (reg_5  ? (~reg_6  & reg_7 ) : (reg_6  & ~reg_7 )) : (reg_5  & (~reg_6  ^ reg_7 )))) | (~reg_1  & ~reg_2  & reg_5  & ~reg_6  & ~reg_7 )) : (reg_5  & ~reg_6  & reg_7  & (~reg_1  | (reg_1  & ~reg_2 )))) : (~reg_6  & ((reg_0  & ~reg_1  & reg_2  & reg_7 ) | (~reg_0  & reg_1  & ~reg_2  & ~reg_7 ) | (~reg_0  & ~reg_1  & reg_2  & ~reg_5  & reg_7 )))) : ((counter_3  & ((reg_0  & ~reg_1  & reg_5  & reg_6  & reg_7 ) | (~reg_0  & reg_1  & ~reg_5  & ~reg_6  & ~reg_7 ))) | (~counter_3  & reg_0  & ~reg_1  & reg_5  & reg_6  & ~reg_7 ) | (reg_1  & ((~reg_7  & (counter_3  ? (reg_2  & (reg_0  ? (reg_5  & ~reg_6 ) : (~reg_5  & reg_6 ))) : (~reg_2  & (reg_0  ? (reg_5  & reg_6 ) : (~reg_5  & ~reg_6 ))))) | (~counter_3  & ~reg_0  & reg_7  & (reg_2  ? (~reg_5  & reg_6 ) : (reg_5  & ~reg_6 ))))) | (counter_3  & ~reg_0  & ~reg_1  & reg_6  & reg_7  & reg_2  & reg_5 )))) | (reg_4  & (reg_0  ? (reg_5  & ((~reg_7  & ((~counter_4  & ((counter_3  & (reg_1  ? (reg_2  & reg_6 ) : (~reg_2  & ~reg_6 ))) | (~counter_3  & ~reg_1  & ~reg_2  & ~reg_6 ))) | (~counter_3  & counter_4  & reg_1  & reg_2  & reg_6 ))) | (counter_3  & counter_4  & reg_7  & (reg_1  ? (~reg_2  & reg_6 ) : (~reg_2  ^ ~reg_6 ))))) : ((reg_7  & (counter_3  ? (~counter_4  & ((~reg_1  & reg_2  & reg_5  & reg_6 ) | (reg_1  & ~reg_2  & ~reg_5  & ~reg_6 ))) : (counter_4  & ((reg_2  & (reg_1  ? (reg_5  & ~reg_6 ) : (~reg_5  & reg_6 ))) | (reg_1  & ~reg_2  & reg_6 ))))) | (~counter_3  & ~reg_7  & ((~reg_2  & ((counter_4  & (reg_1  ? (reg_5  & ~reg_6 ) : (~reg_5  & reg_6 ))) | (~counter_4  & reg_1  & reg_5  & ~reg_6 ))) | (~counter_4  & ~reg_1  & reg_2  & reg_5  & ~reg_6 )))))))) | (~counter_2  & ((counter_4  & (((reg_0  ? (reg_5  & reg_6 ) : (~reg_5  & ~reg_6 )) & ((~counter_3  & ~reg_1  & reg_2  & reg_4  & reg_7 ) | (counter_3  & reg_1  & ~reg_2  & ~reg_4  & ~reg_7 ))) | (reg_2  & (reg_1  ? ((reg_7  & ((reg_0  & ~reg_4  & (counter_3  ? (~reg_5  ^ ~reg_6 ) : (reg_5  & reg_6 ))) | (~counter_3  & ~reg_0  & reg_4  & (~reg_5  ^ reg_6 )))) | (~reg_5  & reg_6  & ~reg_7  & ~counter_3  & ~reg_0  & reg_4 )) : (reg_4  ? ((~reg_7  & ((counter_3  & (reg_0  ? (reg_5  & ~reg_6 ) : (~reg_5  & reg_6 ))) | (~counter_3  & ~reg_0  & reg_5  & ~reg_6 ))) | (~counter_3  & reg_0  & ~reg_5  & reg_7 )) : (~reg_6  & ((counter_3  & (reg_0  ? (reg_5  & ~reg_7 ) : (~reg_5  & reg_7 ))) | (~counter_3  & ~reg_0  & reg_5  & ~reg_7 )))))) | (~reg_2  & (counter_3  ? ((reg_5  & ((reg_4  & ((reg_0  & reg_6  & (~reg_1  ^ reg_7 )) | (~reg_0  & reg_1  & ~reg_6  & reg_7 ))) | (~reg_0  & ~reg_1  & ~reg_4  & reg_6  & reg_7 ))) | (~reg_1  & ~reg_4  & ~reg_5  & (reg_0  ? (~reg_6  & reg_7 ) : (reg_6  & ~reg_7 )))) : ((~reg_5  & ((~reg_1  & ((reg_0  & reg_6  & (~reg_4  ^ reg_7 )) | (~reg_0  & ~reg_4  & ~reg_6  & reg_7 ))) | (~reg_0  & reg_1  & reg_4  & reg_6  & ~reg_7 ))) | (reg_5  & ~reg_6  & ~reg_7  & reg_0  & reg_1  & reg_4 )))))) | (counter_3  & ~counter_4  & ((reg_2  & (reg_5  ? ((~reg_0  & ~reg_1  & ~reg_4  & reg_6  & reg_7 ) | (~reg_6  & ((~reg_1  & (reg_0  ? (~reg_4  ^ reg_7 ) : (reg_4  & ~reg_7 ))) | (~reg_0  & reg_1  & (~reg_4  ^ ~reg_7 ))))) : (reg_6  & ((reg_0  & (reg_1  ? (reg_4  & ~reg_7 ) : (~reg_4  & reg_7 ))) | (~reg_0  & ~reg_1  & reg_4  & reg_7 ))))) | (~reg_0  & ~reg_2  & (((~reg_5  ^ reg_7 ) & (reg_1  ? (~reg_4  & ~reg_6 ) : (reg_4  & reg_6 ))) | (reg_4  & reg_5  & ~reg_7  & (~reg_1  ^ reg_6 )))))))))))) | (~counter_0  & reg_3  & (((~reg_4  ^ ~reg_7 ) & ((reg_0  & ((reg_6  & ((counter_4  & ((counter_2  & (counter_3  ? (reg_1  & ~reg_2 ) : (~reg_1  & reg_2 )) & reg_5 ) | (~counter_2  & ~counter_3  & ~reg_1  & reg_2  & ~reg_5 ))) | (~counter_2  & counter_3  & ~counter_4  & reg_1  & ~reg_2  & reg_5 ))) | (~counter_2  & counter_3  & ~counter_4  & ~reg_1  & ~reg_2  & ~reg_5  & ~reg_6 ))) | (reg_1  & ~reg_2  & ~reg_5  & ~reg_6  & counter_4  & ~reg_0  & counter_2  & counter_3 ))) | (~reg_6  & (counter_2  ? (reg_4  ? ((~reg_2  & (counter_3  ? (counter_4  ? (reg_1  & reg_7  & (reg_0  ^ reg_5 )) : (~reg_1  & ~reg_7  & (~reg_0  ^ reg_5 ))) : ((~reg_0  & ((reg_5  & (counter_4  ? (reg_1  ^ reg_7 ) : (~reg_1  & ~reg_7 ))) | (~counter_4  & reg_1  & ~reg_5  & reg_7 ))) | (counter_4  & reg_0  & reg_1  & ~reg_5  & ~reg_7 )))) | (counter_3  & ~counter_4  & reg_0  & ~reg_1  & reg_2  & ~reg_5  & reg_7 )) : ((reg_5  & (counter_4  ? ((counter_3  & reg_0  & ~reg_1  & reg_2  & reg_7 ) | (~counter_3  & ~reg_0  & reg_1  & ~reg_2  & ~reg_7 )) : ((~reg_0  & ~reg_2  & ~reg_7 ) | (~counter_3  & reg_0  & ~reg_1  & reg_2  & reg_7 )))) | (reg_1  & ~reg_5  & ~reg_7  & ((~counter_3  & ~reg_2  & (~counter_4  ^ reg_0 )) | (counter_3  & counter_4  & ~reg_0  & reg_2 ))))) : (counter_3  ? (reg_2  ? (reg_4  & ((~reg_1  & ((~counter_4  & reg_5  & reg_7 ) | (counter_4  & reg_0  & ~reg_5  & ~reg_7 ))) | (~counter_4  & ~reg_0  & reg_1  & reg_5  & reg_7 ))) : (reg_0  ? ((counter_4  & reg_4  & reg_7  & (reg_1  ^ reg_5 )) | (~counter_4  & reg_1  & ~reg_4  & ~reg_5  & ~reg_7 )) : ((reg_1  & ((reg_4  & (counter_4  ? (reg_5  & ~reg_7 ) : (~reg_5  ^ reg_7 ))) | (counter_4  & ~reg_4  & (~reg_5  ^ ~reg_7 )))) | (counter_4  & ~reg_1  & reg_4  & reg_7 )))) : (counter_4  & (reg_0  ? (((reg_2  ? (reg_4  & ~reg_5 ) : (~reg_4  & reg_5 )) & (~reg_1  ^ reg_7 )) | (~reg_7  & ((~reg_5  & (reg_1  ? (reg_2  ^ reg_4 ) : (~reg_2  & ~reg_4 ))) | (~reg_1  & reg_2  & ~reg_4  & reg_5 )))) : (((~reg_5  ^ ~reg_7 ) & (reg_1  ? (reg_2  & reg_4 ) : (~reg_2  & ~reg_4 ))) | (reg_5  & ((~reg_1  & (reg_2  ? (~reg_4  & reg_7 ) : (reg_4  & ~reg_7 ))) | (reg_1  & ~reg_2  & ~reg_4  & ~reg_7 ))) | (~reg_1  & reg_2  & ~reg_5  & (~reg_4  ^ reg_7 )))))))) | (reg_6  & (reg_0  ? (reg_5  ? (reg_1  ? ((counter_3  & ((~reg_4  & ((counter_2  & reg_2  & reg_7 ) | (~counter_2  & counter_4  & ~reg_2  & ~reg_7 ))) | (~counter_2  & counter_4  & ~reg_2  & reg_4  & ~reg_7 ))) | (~counter_2  & ~counter_3  & counter_4  & reg_2  & ~reg_4  & ~reg_7 )) : (counter_3  ? (reg_2  & ((~counter_2  & counter_4  & (~reg_4  ^ reg_7 )) | (counter_2  & ~counter_4  & reg_4  & reg_7 ))) : ((counter_2  & ~counter_4  & (reg_2  ? (~reg_4  & reg_7 ) : (reg_4  & ~reg_7 ))) | (~counter_2  & counter_4  & ~reg_2  & ~reg_4  & reg_7 )))) : ((counter_3  & ((reg_1  & ((counter_2  & ~reg_7  & (counter_4  ? (~reg_2  & reg_4 ) : (reg_2  & ~reg_4 ))) | (~counter_2  & counter_4  & reg_2  & ~reg_4  & reg_7 ))) | (reg_2  & reg_4  & reg_7  & counter_2  & ~counter_4  & ~reg_1 ))) | (counter_2  & ~counter_3  & ~counter_4  & ~reg_1  & reg_2  & reg_4  & reg_7 ))) : (counter_2  ? (reg_2  ? ((reg_7  & ((counter_4  & ((counter_3  & reg_1  & ~reg_4 ) | (~counter_3  & ~reg_1  & reg_4  & reg_5 ))) | (~counter_3  & ~counter_4  & (reg_1  ? (~reg_4  & reg_5 ) : (reg_4  & ~reg_5 ))))) | (reg_5  & ~reg_7  & ((~counter_4  & ~reg_1  & (counter_3  | (~counter_3  & ~reg_4 ))) | (~counter_3  & counter_4  & reg_1  & ~reg_4 )))) : ((counter_3  & reg_4  & ((~counter_4  & reg_1  & ~reg_5  & reg_7 ) | (~reg_1  & ~reg_5  & reg_7 ) | (reg_1  & reg_5  & ~reg_7 ))) | (~counter_3  & counter_4  & ~reg_1  & ~reg_4  & ~reg_5  & reg_7 ))) : ((counter_4  & ((reg_1  & (counter_3  ? ((reg_2  & ~reg_4  & reg_5  & reg_7 ) | (~reg_2  & reg_4  & ~reg_5  & ~reg_7 )) : (reg_2  ? (reg_4  ? (reg_5  & reg_7 ) : (~reg_5  & ~reg_7 )) : (~reg_4  & reg_7 )))) | (~counter_3  & ~reg_1  & ~reg_4  & (reg_2  ? (~reg_5  & reg_7 ) : (~reg_5  ^ reg_7 ))))) | (reg_2  & ~reg_4  & reg_5  & ~reg_7  & counter_3  & ~counter_4  & reg_1 ))))))))) | (~counter_0  & counter_1  & (reg_4  ? (reg_6  ? (reg_7  ? ((~counter_4  & ((~counter_3  & (counter_2  ? ((reg_0  & ~reg_1  & ~reg_2  & ~reg_3  & reg_5 ) | (~reg_0  & reg_1  & reg_2  & reg_3  & ~reg_5 )) : (~reg_2  & reg_5  & (reg_0  ? (reg_1  & reg_3 ) : (~reg_1  & ~reg_3 ))))) | (~counter_2  & counter_3  & ~reg_2  & ((reg_5  & (reg_0  ? (reg_1  ^ reg_3 ) : (reg_1  & ~reg_3 ))) | (~reg_0  & reg_1  & ~reg_3  & ~reg_5 ))))) | (~counter_2  & counter_4  & ~reg_2  & ((counter_3  & ~reg_0  & (reg_1  ? (~reg_3  & reg_5 ) : (reg_3  & ~reg_5 ))) | (~counter_3  & reg_0  & ~reg_1  & reg_3  & reg_5 )))) : (reg_1  ? (counter_2  ? ((reg_2  & ((counter_3  & ((~counter_4  & reg_0  & ~reg_3  & reg_5 ) | (counter_4  & ~reg_0  & reg_3  & ~reg_5 ))) | (~counter_3  & counter_4  & reg_0  & ~reg_3  & reg_5 ))) | (~counter_3  & ~counter_4  & ~reg_0  & ~reg_2  & ~reg_3  & ~reg_5 )) : ((~reg_2  & ((counter_4  & reg_3  & (counter_3  ? (~reg_0  & reg_5 ) : (reg_0  & ~reg_5 ))) | (~counter_3  & ~counter_4  & ~reg_0  & ~reg_3 ))) | (~counter_3  & ~counter_4  & reg_0  & reg_2  & ~reg_3  & ~reg_5 ))) : ((~counter_2  & ((~reg_2  & ((counter_3  & ~reg_3  & (~counter_4  ^ reg_0 ) & reg_5 ) | (~counter_3  & counter_4  & ~reg_0  & reg_3  & ~reg_5 ))) | (~counter_4  & ~reg_0  & reg_2  & ((reg_3  & (~counter_3  | (counter_3  & reg_5 ))) | (~counter_3  & ~reg_3  & ~reg_5 ))))) | (counter_2  & ~counter_3  & ~counter_4  & ~reg_0  & ~reg_2  & ~reg_3  & reg_5 )))) : ((~reg_2  & (reg_0  ? ((~counter_3  & ((~reg_3  & ((counter_2  & ~reg_1  & reg_5  & reg_7 ) | (~counter_2  & ~counter_4  & reg_1  & ~reg_5  & ~reg_7 ))) | (~counter_2  & ~counter_4  & reg_1  & reg_3  & ~reg_5  & ~reg_7 ))) | (counter_2  & counter_3  & ~reg_1  & ~reg_3  & reg_5  & reg_7 )) : ((reg_1  & (counter_2  ? ((counter_3  & counter_4  & (reg_3  ? (reg_5  & ~reg_7 ) : (~reg_5  & reg_7 ))) | (~counter_3  & ~counter_4  & ~reg_3  & ~reg_5  & reg_7 )) : ((~counter_3  & ~counter_4  & (reg_3  ? (~reg_5  ^ ~reg_7 ) : (~reg_5  ^ reg_7 ))) | (counter_3  & counter_4  & reg_3  & reg_5  & ~reg_7 )))) | (~counter_2  & ~reg_1  & ~reg_3  & reg_5  & reg_7  & (~counter_3  | (counter_3  & counter_4 )))))) | (~counter_2  & ~counter_3  & counter_4  & reg_0  & reg_1  & reg_2  & ~reg_3  & ~reg_5  & ~reg_7 ))) : ((~reg_3  & ((~counter_4  & ((~counter_2  & (reg_0  ? ((~reg_7  & ((~reg_1  & (counter_3  ? (reg_2  ? (~reg_5  & ~reg_6 ) : (reg_5  & reg_6 )) : (reg_2  ? (reg_5  & reg_6 ) : (~reg_5  & ~reg_6 )))) | (~counter_3  & reg_1  & (reg_2  ? (reg_5  & ~reg_6 ) : (~reg_5  & reg_6 ))))) | (~counter_3  & ~reg_2  & reg_6  & reg_7  & (~reg_1  ^ reg_5 ))) : ((~counter_3  & ((~reg_1  & reg_2  & (reg_5  ? (reg_6  & reg_7 ) : (~reg_6  & ~reg_7 ))) | (reg_1  & ~reg_2  & ~reg_5  & ~reg_6  & reg_7 ))) | (counter_3  & ~reg_1  & reg_2  & ~reg_5  & ~reg_6  & reg_7 )))) | (reg_6  & reg_7  & reg_2  & reg_5  & counter_2  & counter_3  & ~reg_0  & ~reg_1 ))) | (~counter_2  & counter_4  & ((~reg_5  & (counter_3  ? (reg_0  & ((~reg_1  & ~reg_6  & (reg_2  ^ reg_7 )) | (reg_1  & ~reg_2  & reg_6  & ~reg_7 ))) : ((~reg_2  & ((reg_0  & reg_6  & reg_7 ) | (~reg_0  & reg_1  & ~reg_6  & ~reg_7 ))) | (~reg_0  & reg_1  & reg_2  & reg_6  & ~reg_7 )))) | (~counter_3  & reg_0  & reg_1  & ~reg_2  & reg_5  & reg_6  & reg_7 ))))) | (~counter_2  & reg_3  & ((~counter_3  & ((~reg_5  & ((counter_4  & reg_2  & ((~reg_0  & ~reg_1  & ~reg_6  & reg_7 ) | (reg_0  & reg_1  & reg_6  & ~reg_7 ))) | (~counter_4  & reg_0  & reg_1  & ~reg_2  & ~reg_6  & ~reg_7 ))) | (reg_2  & reg_5  & reg_6  & (counter_4  ? (reg_0  ? (~reg_1  & reg_7 ) : (reg_1  & ~reg_7 )) : (~reg_0  & ~reg_7 ))))) | (~reg_0  & ~reg_1  & counter_3  & counter_4  & reg_2  & ~reg_5  & ~reg_6  & reg_7 )))))) | (((reg_0  & ~reg_1  & ~reg_2  & ~reg_3  & reg_5 ) | (~reg_0  & reg_1  & reg_2  & reg_3  & ~reg_5 )) & ((~counter_0  & (counter_2  ? ((reg_6  & (counter_1  ? (reg_4  & ((~counter_3  & counter_4  & reg_7  & reg_8 ) | (counter_3  & ~counter_4  & ~reg_7  & ~reg_8 ))) : (counter_4  & ~reg_4  & (counter_3  ? (~reg_7  & ~reg_8 ) : (reg_7  & reg_8 ))))) | (~counter_1  & counter_3  & ~reg_6  & (counter_4  ? (reg_4  ? (~reg_7  & ~reg_8 ) : (reg_7  & reg_8 )) : (~reg_4  & (~reg_7  ^ reg_8 ))))) : ((reg_6  & reg_7  & reg_8  & (counter_1  ? (counter_3  ? (counter_4  & reg_4 ) : (~counter_4  & ~reg_4 )) : (counter_3  ? (~counter_4  & ~reg_4 ) : (counter_4  & reg_4 )))) | (~counter_1  & ~counter_3  & counter_4  & reg_4  & ~reg_6  & ~reg_7  & ~reg_8 )))) | (counter_0  & ~counter_1  & ~counter_2  & ~counter_3  & ~counter_4  & reg_4  & reg_6  & ~reg_7  & ~reg_8 ))) | (~counter_0  & (counter_2  ? ((~counter_3  & (reg_2  ? ((~reg_3  & ((reg_5  & ((reg_7  & reg_8  & (counter_1  ? ((~reg_0  & ~reg_1  & ~reg_4  & reg_6 ) | (reg_0  & reg_1  & reg_4  & ~reg_6 )) : ((reg_1  & ((~reg_0  & reg_4  & reg_6 ) | (~reg_6  & (reg_0  | (~reg_0  & ~reg_4 ))))) | (reg_0  & ~reg_1  & reg_4  & ~reg_6 )))) | (~counter_1  & ~reg_7  & ~reg_8  & (reg_0  ? (reg_1  ? (~reg_4  & ~reg_6 ) : (reg_4  & reg_6 )) : (reg_1  & ~reg_6 ))))) | (~counter_1  & ~reg_5  & ((reg_0  & ((reg_6  & ((reg_1  & reg_7  & (reg_4  ^ reg_8 )) | (~reg_7  & ~reg_8  & ~reg_1  & reg_4 ))) | (~reg_1  & reg_4  & ~reg_6  & (~reg_7  ^ reg_8 )))) | (~reg_0  & reg_1  & reg_4  & reg_6  & reg_7  & reg_8 ))))) | (~counter_1  & reg_3  & ((~reg_6  & (((reg_0  ^ reg_5 ) & ((~reg_7  & ~reg_8  & ~reg_1  & reg_4 ) | (reg_1  & ~reg_4  & reg_7  & reg_8 ))) | (reg_0  & reg_1  & (reg_4  ^ reg_5 ) & (~reg_7  ^ reg_8 )))) | (reg_0  & ~reg_4  & reg_6  & ((reg_1  & (~reg_7  ^ reg_8 )) | (~reg_1  & ~reg_5  & ~reg_7  & ~reg_8 )))))) : ((~reg_5  & ((~reg_1  & (((reg_6  ? (~reg_7  & ~reg_8 ) : (reg_7  & reg_8 )) & ((~counter_1  & reg_3  & (reg_0  ^ reg_4 )) | (~reg_3  & reg_4  & counter_1  & reg_0 ))) | (~counter_1  & ((reg_3  & ((~reg_0  & reg_6  & (reg_4  ? (reg_7  & reg_8 ) : (~reg_7  & ~reg_8 ))) | (reg_0  & ~reg_4  & ~reg_6  & ~reg_7  & ~reg_8 ))) | (reg_0  & ~reg_3  & reg_4  & (reg_6  ? (reg_7  & reg_8 ) : (~reg_7  & ~reg_8 ))))) | (counter_1  & reg_0  & reg_3  & ~reg_4  & ~reg_6  & ~reg_7  & ~reg_8 ))) | (~counter_1  & reg_1  & ((~reg_4  & ((reg_7  & reg_8  & (reg_0  ? ~reg_6  : (reg_3  & reg_6 ))) | (~reg_0  & reg_3  & reg_6  & ~reg_7  & ~reg_8 ))) | (reg_6  & ~reg_7  & ~reg_8  & reg_0  & ~reg_3  & reg_4 ))))) | (~counter_1  & reg_5  & ((reg_7  & reg_8  & ((reg_0  & reg_3  & ~reg_6  & (~reg_1  ^ ~reg_4 )) | (~reg_0  & reg_1  & ~reg_3  & ~reg_4  & reg_6 ))) | (reg_0  & ~reg_1  & reg_3  & reg_4  & ~reg_6  & ~reg_7  & ~reg_8 )))))) | (~counter_1  & counter_3  & (reg_3  ? ((~reg_6  & ((reg_2  & ((~reg_7  & ~reg_8  & ((reg_0  & reg_1  & ~reg_4 ) | (~reg_0  & ~reg_1  & reg_4  & ~reg_5 ))) | (~reg_0  & ~reg_1  & reg_4  & reg_5  & reg_7  & reg_8 ))) | (reg_0  & ~reg_2  & ~reg_4  & ~reg_7  & ~reg_8  & (~reg_1  ^ reg_5 )))) | (reg_1  & reg_6  & ((~reg_0  & reg_7  & reg_8  & (reg_2  ? (reg_4  & reg_5 ) : (~reg_4  & ~reg_5 ))) | (reg_0  & ~reg_2  & ~reg_4  & reg_5  & ~reg_7  & ~reg_8 )))) : (reg_2  ? (((reg_0  ^ reg_4 ) & ((~reg_1  & ~reg_5  & ~reg_6  & reg_7  & reg_8 ) | (reg_1  & reg_5  & reg_6  & ~reg_7  & ~reg_8 ))) | (~reg_0  & ((reg_4  & ((reg_1  & reg_5  & ~reg_6  & reg_7  & reg_8 ) | (~reg_1  & ~reg_5  & reg_6  & ~reg_7  & ~reg_8 ))) | (reg_1  & ~reg_4  & reg_5  & ~reg_6  & (~reg_7  ^ reg_8 ))))) : ((~reg_5  & ((reg_4  & (reg_0  ? (~reg_1  & (reg_6  ? (~reg_7  & ~reg_8 ) : (reg_7  & reg_8 ))) : (reg_1  & (reg_6  ? (reg_7  & reg_8 ) : (~reg_7  & ~reg_8 ))))) | (~reg_0  & reg_1  & ~reg_4  & reg_6  & (~reg_7  ^ reg_8 )))) | (~reg_0  & ~reg_4  & reg_5  & reg_6  & (reg_1  ? (~reg_7  ^ reg_8 ) : (~reg_7  & ~reg_8 )))))))) : (((reg_6  ? (~reg_7  & ~reg_8 ) : (reg_7  & reg_8 )) & ((counter_3  & ((~counter_1  & ~reg_4  & ((~reg_0  & ~reg_1  & ~reg_2  & reg_3  & reg_5 ) | (reg_0  & reg_1  & reg_2  & ~reg_3  & ~reg_5 ))) | (counter_1  & reg_0  & ~reg_1  & ~reg_2  & ~reg_3  & reg_4  & ~reg_5 ))) | (counter_1  & ~counter_3  & ~reg_1  & ~reg_3  & reg_5  & (reg_0  ? (~reg_2  & reg_4 ) : (reg_2  & ~reg_4 ))))) | (reg_3  & (reg_1  ? (counter_1  ? (reg_0  ? (~reg_4  & ((~counter_3  & reg_7  & reg_8  & (reg_2  ? (~reg_5  & reg_6 ) : (reg_5  & ~reg_6 ))) | (~reg_6  & ~reg_7  & ~reg_8  & counter_3  & ~reg_2  & reg_5 ))) : ((reg_4  & ((reg_2  & reg_5  & ((counter_3  & ~reg_6  & (~reg_7  ^ reg_8 )) | (~reg_7  & ~reg_8  & ~counter_3  & reg_6 ))) | (reg_6  & reg_7  & reg_8  & ~counter_3  & ~reg_2  & ~reg_5 ))) | (~counter_3  & ~reg_2  & ~reg_4  & ~reg_5  & ~reg_6  & ~reg_7  & ~reg_8 ))) : (counter_3  & ((~reg_6  & ((~reg_5  & ((reg_4  & ((reg_0  & (reg_2  ? (reg_7  & reg_8 ) : (~reg_7  & ~reg_8 ))) | (~reg_0  & reg_2  & ~reg_7  & ~reg_8 ))) | (~reg_0  & ~reg_2  & ~reg_4  & ~reg_7  & ~reg_8 ))) | (reg_5  & ~reg_7  & ~reg_8  & reg_0  & reg_2  & ~reg_4 ))) | (~reg_0  & ~reg_2  & reg_6  & ((~reg_4  & (reg_5  ? (reg_7  & reg_8 ) : (~reg_7  & ~reg_8 ))) | (reg_4  & reg_5  & reg_7  & reg_8 )))))) : ((~reg_5  & ((reg_7  & reg_8  & ((reg_0  & ((~reg_2  & ((counter_1  & ~reg_4  & ~reg_6 ) | (~counter_1  & counter_3  & reg_4  & reg_6 ))) | (~counter_1  & counter_3  & reg_2  & ~reg_4  & reg_6 ))) | (counter_1  & ~counter_3  & ~reg_0  & reg_2  & reg_4  & ~reg_6 ))) | (~reg_2  & ~reg_4  & ~reg_7  & ~reg_8  & ((~reg_6  & (counter_1  ? (~counter_3  ^ reg_0 ) : (counter_3  & ~reg_0 ))) | (~counter_1  & counter_3  & reg_0  & reg_6 ))))) | (~counter_1  & counter_3  & reg_5  & ((reg_6  & ((~reg_7  & ~reg_8  & (reg_0  ? ~reg_2  : (reg_2  & reg_4 ))) | (~reg_0  & reg_2  & reg_4  & reg_7  & reg_8 ))) | (~reg_6  & ~reg_7  & ~reg_8  & ~reg_0  & ~reg_2  & reg_4 )))))) | (~reg_3  & (reg_5  ? ((~reg_7  & ~reg_8  & ((reg_0  & ~reg_1  & ((counter_1  & ~counter_3  & ~reg_2  & (reg_4  ^ reg_6 )) | (~counter_1  & counter_3  & reg_2  & reg_4  & reg_6 ))) | (~counter_1  & counter_3  & ~reg_0  & reg_1  & reg_4  & (~reg_2  ^ reg_6 )))) | (counter_3  & reg_1  & reg_2  & reg_6  & reg_7  & reg_8  & (counter_1  ? (reg_0  & ~reg_4 ) : (~reg_0  & reg_4 )))) : (reg_2  ? ((reg_0  & ((~reg_1  & ((~counter_1  & counter_3  & reg_7  & reg_8  & (~reg_4  ^ reg_6 )) | (~reg_6  & ~reg_7  & ~reg_8  & counter_1  & ~counter_3  & ~reg_4 ))) | (counter_1  & ~counter_3  & reg_1  & ((~reg_4  & ~reg_6  & ~reg_7  & ~reg_8 ) | (reg_4  & reg_6  & reg_7  & reg_8 ))))) | (counter_3  & ~reg_0  & ((~reg_7  & ~reg_8  & ((~counter_1  & ~reg_4  & reg_6 ) | (reg_4  & ~reg_6  & counter_1  & ~reg_1 ))) | (~counter_1  & reg_1  & reg_7  & reg_8  & (reg_4  ^ reg_6 ))))) : ((reg_4  & ((counter_3  & (reg_0  ? (reg_6  & ((reg_7  & reg_8  & counter_1  & ~reg_1 ) | (~reg_7  & ~reg_8  & ~counter_1  & reg_1 ))) : (~reg_6  & (~reg_7  ^ reg_8 ) & (counter_1  ^ ~reg_1 )))) | (counter_1  & ~counter_3  & reg_0  & reg_7  & reg_8  & ~reg_1  & reg_6 ))) | (~reg_4  & ~reg_6  & ~reg_7  & ~reg_8  & reg_0  & reg_1  & ~counter_1  & counter_3 )))))))) | (~counter_3  & ~reg_0  & reg_1  & counter_0  & ~counter_1  & ~counter_2  & reg_2  & reg_3  & reg_4  & ~reg_5  & ~reg_6  & reg_7  & reg_8 ) | (~counter_0  & (counter_4  ? (reg_4  ? (counter_3  ? (counter_2  ? (counter_1  ? ((~reg_5  & ~reg_6  & reg_7  & reg_8  & ~reg_0  & reg_1  & reg_2  & reg_3 ) | (reg_0  & ~reg_1  & ~reg_2  & ~reg_3  & reg_5  & reg_6  & ~reg_7  & ~reg_8 )) : (reg_2  ? (reg_1  ? ((~reg_3  & (((reg_6  ? (reg_7  & reg_8 ) : (~reg_7  & ~reg_8 )) & (~reg_0  | (reg_0  & reg_5 ))) | (~reg_0  & ~reg_5  & reg_6  & ~reg_7  & ~reg_8 ))) | (reg_6  & ~reg_7  & ~reg_8  & ~reg_0  & reg_3  & reg_5 )) : (reg_0  ? ((~reg_5  & ((~reg_7  & (reg_3  ? reg_8  : (reg_6  & ~reg_8 ))) | (~reg_3  & ~reg_6  & reg_7  & reg_8 ))) | (reg_3  & reg_5  & (reg_6  ? (~reg_7  & reg_8 ) : (~reg_7  ^ reg_8 )))) : (reg_6  & ((~reg_7  & (reg_3  ? ~reg_8  : (reg_5  & reg_8 ))) | (reg_7  & ~reg_8  & reg_3  & ~reg_5 ))))) : (reg_7  ? ((reg_3  & ((reg_6  & ((reg_8  & (reg_0  ? (reg_1  ^ reg_5 ) : (reg_1  & reg_5 ))) | (~reg_0  & reg_1  & ~reg_5  & ~reg_8 ))) | (~reg_0  & ~reg_1  & ~reg_6  & (reg_5  ^ ~reg_8 )))) | (~reg_1  & ~reg_3  & reg_8  & (reg_0  ? (~reg_5  ^ ~reg_6 ) : (reg_5  & reg_6 )))) : ((reg_1  & ((~reg_8  & ((~reg_0  & ~reg_5  & reg_6 ) | (~reg_6  & (reg_0  ? (reg_3  | (~reg_3  & ~reg_5 )) : (~reg_3  & reg_5 ))))) | (reg_0  & ~reg_3  & reg_5  & ~reg_6  & reg_8 ))) | (~reg_0  & ~reg_1  & reg_3  & reg_5  & reg_6  & ~reg_8 ))))) : (reg_0  ? (reg_2  ? ((~counter_1  & ((~reg_5  & ((~reg_6  & ((reg_1  & ~reg_7  & (~reg_3  ^ ~reg_8 )) | (~reg_1  & reg_3  & reg_7  & reg_8 ))) | (~reg_1  & reg_3  & reg_6  & ~reg_7  & ~reg_8 ))) | (reg_1  & ~reg_3  & reg_5  & reg_7  & (reg_6  ^ reg_8 )))) | (reg_5  & reg_6  & ~reg_7  & ~reg_8  & counter_1  & reg_1  & ~reg_3 )) : ((reg_3  & (((counter_1  ^ ~reg_1 ) & ((~reg_5  & ~reg_6  & ~reg_7  & ~reg_8 ) | (reg_5  & reg_6  & reg_7  & reg_8 ))) | (~reg_1  & ((~counter_1  & ~reg_5  & (reg_6  ? (~reg_7  & ~reg_8 ) : (reg_7  & reg_8 ))) | (reg_6  & reg_7  & reg_8  & counter_1  & reg_5 ))))) | (~counter_1  & reg_1  & ~reg_3  & ((~reg_5  & reg_7  & reg_8 ) | (reg_5  & ~reg_6  & ~reg_7  & ~reg_8 ))))) : (reg_1  ? ((~reg_5  & ((reg_6  & ((~reg_2  & ((counter_1  & (reg_3  ? (reg_7  & ~reg_8 ) : (~reg_7  & reg_8 ))) | (reg_7  & reg_8  & ~counter_1  & reg_3 ))) | (~counter_1  & reg_2  & ~reg_3  & ~reg_8 ))) | (reg_2  & ~reg_3  & ~reg_6  & ~reg_7  & ~reg_8 ))) | (~counter_1  & ~reg_2  & ~reg_3  & reg_5  & reg_6  & (~reg_7  ^ reg_8 ))) : ((reg_7  & (counter_1  ? ((reg_2  & reg_3  & ~reg_5  & ~reg_6  & reg_8 ) | (~reg_2  & ~reg_3  & reg_5  & reg_6  & ~reg_8 )) : (reg_8  & ((reg_2  & (reg_5  ? (reg_3  ^ reg_6 ) : reg_3 )) | (~reg_2  & reg_3  & ~reg_5  & reg_6 ))))) | (~counter_1  & ~reg_7  & ((reg_6  & ((~reg_2  & reg_3  & ~reg_8 ) | (reg_2  & ~reg_3  & reg_5  & reg_8 ))) | (reg_2  & ~reg_3  & ~reg_6  & (reg_5  ^ ~reg_8 )))))))) : (reg_2  ? ((~counter_2  & (reg_5  ? (reg_0  ? ((~reg_3  & ((reg_1  & ((~reg_8  & (counter_1  ? (~reg_6  ^ reg_7 ) : (~reg_6  & reg_7 ))) | (reg_7  & reg_8  & ~counter_1  & reg_6 ))) | (~counter_1  & ~reg_1  & (reg_6  ? (~reg_7  & ~reg_8 ) : (reg_7  & reg_8 ))))) | (~counter_1  & ~reg_1  & reg_3  & (reg_6  ? (~reg_7  & ~reg_8 ) : reg_8 ))) : ((~reg_6  & ((reg_8  & ((reg_3  & ((reg_7  & (counter_1  | (~counter_1  & reg_1 ))) | (~counter_1  & ~reg_1  & ~reg_7 ))) | (counter_1  & reg_1  & ~reg_3  & reg_7 ))) | (~counter_1  & reg_1  & ~reg_3  & ~reg_7  & ~reg_8 ))) | (~counter_1  & reg_6  & ~reg_7  & (reg_1  ? (reg_3  & ~reg_8 ) : (~reg_3  ^ reg_8 ))))) : ((~reg_7  & ~reg_8  & ((~reg_0  & ((~reg_6  & (counter_1  ? (reg_1  ^ reg_3 ) : (~reg_1  & ~reg_3 ))) | (~counter_1  & reg_3  & reg_6 ))) | (~counter_1  & reg_0  & reg_1  & ~reg_6 ))) | (~counter_1  & ~reg_1  & reg_3  & reg_6  & reg_7  & reg_8 )))) | (~counter_1  & counter_2  & ((reg_6  & ((reg_8  & ((reg_7  & ((reg_0  & ~reg_3  & (~reg_1  ^ reg_5 )) | (~reg_0  & reg_1  & reg_3  & reg_5 ))) | (reg_0  & ~reg_1  & reg_3  & ~reg_5  & ~reg_7 ))) | (~reg_0  & reg_1  & ~reg_3  & ~reg_7  & ~reg_8 ))) | (~reg_0  & ~reg_1  & reg_5  & ~reg_6  & (reg_3  ? (reg_7  & reg_8 ) : ~reg_8 ))))) : (reg_5  ? (reg_6  ? ((((~reg_7  & ((~counter_2  & (reg_0  ? (reg_1  & reg_8 ) : (~reg_1  & ~reg_8 ))) | (counter_2  & reg_0  & ~reg_1  & ~reg_8 ))) | (~counter_2  & ~reg_0  & reg_1  & reg_7  & reg_8 )) & (counter_1  ^ reg_3 )) | (reg_7  & ((reg_1  & ((~counter_2  & (counter_1  ? (reg_3  & (~reg_0  ^ reg_8 )) : (~reg_3  & reg_8 ))) | (~counter_1  & counter_2  & ~reg_0  & reg_3  & ~reg_8 ))) | (~counter_1  & counter_2  & ~reg_1  & reg_8  & (reg_0  | (~reg_0  & reg_3 ))))) | (~counter_1  & counter_2  & ~reg_7  & ~reg_8  & (reg_0  ? reg_1  : (~reg_1  & reg_3 )))) : ((~counter_1  & (reg_1  ? ((reg_3  & (counter_2  ? (reg_0  ? (~reg_7  & ~reg_8 ) : (reg_7  & reg_8 )) : (reg_7  & (reg_0  ^ reg_8 )))) | (~counter_2  & ~reg_3  & (reg_0  ? (reg_7  & reg_8 ) : (~reg_7  ^ reg_8 )))) : ((~reg_0  & ((~reg_7  & ~reg_8  & (counter_2  | (~counter_2  & ~reg_3 ))) | (reg_7  & reg_8  & ~counter_2  & ~reg_3 ))) | (~counter_2  & reg_0  & ~reg_3  & reg_7  & reg_8 )))) | (counter_1  & ~counter_2  & ~reg_0  & reg_1  & reg_3  & reg_7  & ~reg_8 ))) : (reg_0  ? (((reg_6  ? (~reg_7  & ~reg_8 ) : (reg_7  & reg_8 )) & ((~counter_1  & (counter_2  ? (~reg_1  & reg_3 ) : (reg_1  & ~reg_3 ))) | (counter_1  & ~counter_2  & ~reg_1  & ~reg_3 ))) | (~counter_1  & (((~reg_3  ^ reg_6 ) & ((counter_2  & reg_1  & reg_7  & reg_8 ) | (~counter_2  & ~reg_1  & ~reg_7  & ~reg_8 ))) | (~counter_2  & (reg_3  ? ((reg_7  & (reg_1  ? reg_8  : (reg_6  & ~reg_8 ))) | (~reg_7  & reg_8  & ~reg_1  & ~reg_6 )) : (~reg_8  & (reg_1  ? (~reg_6  ^ reg_7 ) : (reg_6  & ~reg_7 ))))))) | (counter_1  & ~counter_2  & reg_1  & ~reg_3  & ~reg_6  & ~reg_7  & ~reg_8 )) : (reg_1  ? (reg_6  ? ((~counter_2  & ((~reg_3  & (counter_1  ? (~reg_7  ^ reg_8 ) : (reg_7  & reg_8 ))) | (~reg_7  & ~reg_8  & ~counter_1  & reg_3 ))) | (counter_1  & counter_2  & (reg_3  ? (reg_7  & reg_8 ) : (~reg_7  & ~reg_8 )))) : ((reg_8  & ((~reg_3  & (counter_1  ? (counter_2  ^ reg_7 ) : reg_7 )) | (~counter_1  & ~counter_2  & reg_3 ))) | (~counter_1  & counter_2  & ~reg_3  & ~reg_7  & ~reg_8 ))) : ((~counter_1  & ((~counter_2  & (reg_7  ? (reg_3  ? (reg_6  & reg_8 ) : (~reg_6  & ~reg_8 )) : ((~reg_8  & (reg_3  | (~reg_3  & ~reg_6 ))) | (~reg_3  & reg_6  & reg_8 )))) | (counter_2  & ~reg_3  & reg_6  & reg_7  & reg_8 ))) | (~reg_6  & reg_7  & reg_8  & counter_1  & ~counter_2  & reg_3 ))))))) : (counter_2  ? ((~counter_1  & (counter_3  ? (reg_2  ? (reg_7  ? ((reg_3  & (reg_0  ? (~reg_5  & (reg_1  ? (reg_6  ^ reg_8 ) : (~reg_6  & reg_8 ))) : (reg_5  & (reg_1  ? (~reg_6  & reg_8 ) : (reg_6  & ~reg_8 ))))) | (reg_1  & ~reg_3  & ((~reg_5  & (~reg_0  ^ reg_8 )) | (~reg_0  & reg_5  & reg_6  & reg_8 )))) : ((~reg_8  & ((~reg_6  & ((~reg_0  & reg_1  & reg_3  & reg_5 ) | (~reg_1  & (reg_0  ? (~reg_3  ^ reg_5 ) : (~reg_3  & ~reg_5 ))))) | (~reg_1  & ~reg_3  & reg_6  & (~reg_0  ^ reg_5 )))) | (~reg_0  & ~reg_1  & ~reg_3  & reg_5  & reg_6  & reg_8 ))) : ((~reg_8  & (reg_0  ? (~reg_3  & ~reg_5  & (reg_1  ? (reg_6  & reg_7 ) : ~reg_7 )) : ((reg_3  & (reg_1  ? (reg_5  & ~reg_6 ) : (~reg_5  & reg_6 ))) | (reg_1  & ~reg_3  & ~reg_5  & ~reg_6  & ~reg_7 )))) | (reg_7  & reg_8  & ((~reg_1  & reg_6  & (reg_0  ? ~reg_3  : (reg_3  & reg_5 ))) | (~reg_0  & reg_1  & ~reg_3  & ~reg_5  & ~reg_6 ))))) : (reg_6  ? (reg_3  ? (reg_0  ? (reg_1  & ~reg_2  & ((~reg_5  & ~reg_7  & ~reg_8 ) | (reg_8  & (reg_5  | (~reg_5  & reg_7 ))))) : (reg_2  & ((~reg_7  & reg_8  & reg_1  & ~reg_5 ) | (reg_7  & ~reg_8  & ~reg_1  & reg_5 )))) : (reg_8  & (reg_1  ? (reg_2  & (reg_0  ? (~reg_5  ^ reg_7 ) : reg_7 )) : (reg_2  ? reg_7  : (reg_0  ? (~reg_5  & reg_7 ) : (reg_5  & ~reg_7 )))))) : (reg_1  ? ((~reg_3  & ((~reg_0  & reg_2  & ~reg_5  & reg_7  & reg_8 ) | (reg_0  & ~reg_2  & reg_5  & ~reg_7  & ~reg_8 ))) | (~reg_0  & reg_3  & ((~reg_8  & (reg_2  ? (~reg_5  ^ ~reg_7 ) : (~reg_5  & ~reg_7 ))) | (reg_7  & reg_8  & ~reg_2  & ~reg_5 )))) : (reg_0  ? ((~reg_2  & reg_5  & reg_7  & reg_8 ) | (reg_2  & ~reg_5  & ~reg_7  & ~reg_8 ) | (~reg_2  & ~reg_3  & ~reg_5  & ~reg_7  & reg_8 )) : (((reg_2  ^ reg_7 ) & (reg_3  ? (~reg_5  & reg_8 ) : (reg_5  & ~reg_8 ))) | (reg_5  & ~reg_8  & (reg_2  ? (~reg_3  & reg_7 ) : (reg_3  & ~reg_7 ))))))))) | (reg_0  & reg_1  & ~reg_2  & counter_1  & ~counter_3  & reg_3  & ~reg_5  & reg_6  & reg_7  & reg_8 )) : (reg_7  ? ((reg_8  & ((((reg_1  & ~reg_2  & reg_5  & reg_6 ) | (~reg_1  & reg_2  & ~reg_5  & ~reg_6 )) & ((counter_1  & (counter_3  ? (reg_0  & reg_3 ) : (~reg_0  & ~reg_3 ))) | (reg_0  & reg_3  & ~counter_1  & counter_3 ))) | (~counter_3  & (((reg_1  ? (reg_3  & reg_6 ) : (~reg_3  & ~reg_6 )) & ((counter_1  & ~reg_2  & (reg_0  ^ reg_5 )) | (reg_2  & reg_5  & ~counter_1  & reg_0 ))) | (~counter_1  & ((~reg_1  & (reg_0  ? (reg_2  ? (reg_5  & reg_6 ) : (~reg_5  & ~reg_6 )) : (reg_2  & (~reg_5  ^ reg_6 )))) | (~reg_0  & reg_1  & ~reg_2  & ~reg_5  & ~reg_6 ) | (~reg_3  & ((reg_1  & ((reg_5  & ~reg_6 ) | (reg_0  & ~reg_2  & ~reg_5  & reg_6 ))) | (reg_0  & ~reg_1  & (reg_2  ? (~reg_5  & ~reg_6 ) : reg_6 )))) | (reg_0  & ~reg_1  & reg_2  & reg_3  & reg_5  & ~reg_6 ))) | (reg_2  & ~reg_3  & reg_5  & reg_6  & counter_1  & ~reg_0  & reg_1 ))) | (~counter_1  & counter_3  & ((~reg_6  & (((~reg_1  ^ reg_2 ) & (reg_0  ? (reg_3  & ~reg_5 ) : (~reg_3  & reg_5 ))) | (~reg_0  & reg_2  & (reg_1  ? (reg_3  & ~reg_5 ) : (~reg_3  & reg_5 ))))) | (reg_0  & reg_6  & ((~reg_1  & (reg_2  ? (~reg_3  & ~reg_5 ) : reg_3 )) | (reg_1  & ~reg_2  & reg_3  & ~reg_5 ))))))) | (~counter_1  & ~reg_8  & (counter_3  ? ((reg_0  & ((~reg_2  & ((reg_1  & ~reg_6  & (~reg_3  ^ ~reg_5 )) | (~reg_1  & ~reg_3  & reg_5  & reg_6 ))) | (~reg_1  & reg_2  & ~reg_3  & reg_5  & reg_6 ))) | (~reg_0  & ~reg_1  & reg_2  & reg_3  & reg_5  & reg_6 )) : ((reg_2  & ((reg_1  & ~reg_6  & (reg_0  ? (~reg_3  ^ reg_5 ) : (reg_3  & reg_5 ))) | (~reg_0  & ~reg_1  & ~reg_3  & ~reg_5  & reg_6 ))) | (reg_0  & ~reg_2  & reg_3  & ~reg_5  & reg_6 ))))) : (reg_5  ? (counter_3  ? ((~counter_1  & (reg_0  ? ((reg_3  & ((~reg_1  & ~reg_6  & ~reg_8 ) | (reg_1  & reg_2  & reg_6  & reg_8 ))) | (~reg_1  & ~reg_2  & ~reg_3  & ~reg_6  & reg_8 )) : ((~reg_3  & (reg_1  ? (reg_2  ? (~reg_6  & ~reg_8 ) : (reg_6  ^ reg_8 )) : (reg_2  ? (~reg_6  & reg_8 ) : (reg_6  & ~reg_8 )))) | (reg_1  & ~reg_2  & reg_3  & reg_6  & ~reg_8 )))) | (counter_1  & ~reg_0  & ~reg_1  & reg_2  & ~reg_3  & reg_6  & reg_8 )) : (reg_1  ? ((reg_0  & ((reg_3  & ((counter_1  & (reg_2  ? (~reg_6  & ~reg_8 ) : (reg_6  & reg_8 ))) | (~counter_1  & ~reg_2  & reg_6  & ~reg_8 ))) | (~counter_1  & ~reg_3  & (reg_2  ? (~reg_6  & reg_8 ) : (~reg_6  ^ reg_8 ))))) | (~counter_1  & ~reg_0  & ((~reg_3  & ((reg_8  & (reg_2  | (~reg_2  & reg_6 ))) | (~reg_2  & ~reg_6  & ~reg_8 ))) | (reg_2  & reg_3  & ~reg_6  & ~reg_8 )))) : ((~counter_1  & (reg_0  ? ((reg_2  & (reg_3  ? (reg_6  & ~reg_8 ) : (~reg_6  & reg_8 ))) | (~reg_2  & ~reg_3  & ~reg_6  & ~reg_8 )) : (~reg_2  & ~reg_8  & (~reg_3  | (reg_3  & reg_6 ))))) | (counter_1  & ~reg_0  & ~reg_2  & ~reg_3  & reg_6  & ~reg_8 )))) : ((~reg_8  & (reg_6  ? ((~counter_1  & (counter_3  ? ((reg_0  & ~reg_1  & ~reg_2  & ~reg_3 ) | (~reg_0  & reg_1  & reg_2  & reg_3 )) : (reg_0  ? (reg_1  ? (reg_2  & ~reg_3 ) : (~reg_2  & reg_3 )) : (reg_1  ? (~reg_2  & ~reg_3 ) : (reg_2  & reg_3 ))))) | (reg_1  & ~reg_2  & reg_3  & counter_1  & ~counter_3  & reg_0 )) : (counter_3  ? (counter_1  ? ((reg_0  & reg_1  & reg_2  & ~reg_3 ) | (~reg_0  & ~reg_1  & ~reg_2  & reg_3 )) : (reg_2  & (reg_0  ? (~reg_1  & ~reg_3 ) : (~reg_1  | (reg_1  & ~reg_3 ))))) : ((reg_0  & ((counter_1  & ~reg_1  & reg_3 ) | (~counter_1  & reg_1  & ~reg_3 ) | (~reg_1  & ~reg_3  & (counter_1  ^ reg_2 )))) | (~counter_1  & ~reg_0  & reg_1  & ~reg_2  & reg_3 ))))) | (~counter_1  & ~counter_3  & reg_8  & ((reg_2  & ((reg_1  & (reg_0  ? (reg_3  & reg_6 ) : ~reg_3 )) | (reg_0  & ~reg_1  & (reg_3  ^ reg_6 )))) | (~reg_0  & reg_1  & ~reg_2  & ~reg_3  & ~reg_6 )))))))) : (counter_3  ? (reg_5  ? (reg_0  ? (reg_2  ? (((~reg_7  ^ reg_8 ) & ((~reg_6  & ((~counter_2  & ((counter_1  & (reg_1  ^ reg_3 ) & reg_4 ) | (~counter_1  & reg_1  & ~reg_3  & ~reg_4 ))) | (~counter_1  & counter_2  & ~reg_1  & ~reg_3  & ~reg_4 ))) | (~counter_1  & counter_2  & ~reg_1  & reg_3  & ~reg_4  & reg_6 ))) | (~counter_1  & (reg_3  ? ((~reg_4  & ((~reg_7  & (counter_2  ? (reg_1  ? (reg_6  & ~reg_8 ) : (~reg_6  & reg_8 )) : (~reg_1  & reg_8 ))) | (counter_2  & reg_1  & ~reg_6  & reg_7  & reg_8 ))) | (~reg_1  & reg_4  & reg_6  & (counter_2  ? (~reg_7  & ~reg_8 ) : (reg_7  & reg_8 )))) : ((reg_4  & ((counter_2  & ~reg_1  & reg_7  & reg_8 ) | (~counter_2  & reg_1  & ~reg_7  & ~reg_8 ) | (~counter_2  & ~reg_1  & ~reg_6  & ~reg_7  & ~reg_8 ))) | (reg_6  & reg_7  & reg_8  & ~counter_2  & ~reg_1  & ~reg_4 )))) | (~reg_4  & ~reg_6  & ~reg_7  & ~reg_8  & counter_1  & ~counter_2  & reg_1  & reg_3 )) : (counter_1  ? (counter_2  ? ((reg_6  & reg_7  & reg_8  & ~reg_1  & ~reg_3  & reg_4 ) | (~reg_6  & ~reg_7  & ~reg_8  & reg_1  & reg_3  & ~reg_4 )) : ((reg_6  & ((~reg_3  & ((reg_1  & ~reg_4  & reg_7  & reg_8 ) | (~reg_1  & reg_4  & (~reg_7  ^ reg_8 )))) | (reg_1  & reg_3  & ~reg_4  & ~reg_8 ))) | (~reg_1  & ~reg_3  & reg_4  & ~reg_6  & (~reg_7  ^ reg_8 )))) : ((((reg_1  & reg_7  & (~reg_3  ^ reg_4 )) | (~reg_1  & reg_3  & ~reg_4  & ~reg_7 )) & (counter_2  ? (reg_6  & ~reg_8 ) : (~reg_6  & reg_8 ))) | (reg_4  & (counter_2  ? ((~reg_1  & reg_3  & reg_6  & ~reg_7  & ~reg_8 ) | (reg_8  & ((reg_1  & (reg_3  ? (~reg_6  & reg_7 ) : (reg_6  & ~reg_7 ))) | (~reg_1  & ~reg_3  & reg_6  & reg_7 )))) : ((~reg_6  & (reg_1  ? (reg_3  ? (~reg_7  & ~reg_8 ) : (reg_7  & reg_8 )) : (reg_8  & (~reg_3  ^ reg_7 )))) | (~reg_3  & reg_6  & reg_7  & (~reg_1  ^ reg_8 ))))) | (~counter_2  & ~reg_4  & ((~reg_6  & ((reg_3  & (reg_1  ? (~reg_7  ^ reg_8 ) : (reg_7  & reg_8 ))) | (~reg_1  & ~reg_3  & reg_7  & ~reg_8 ))) | (reg_1  & reg_6  & (reg_3  ? (~reg_7  & ~reg_8 ) : (reg_7  & reg_8 )))))))) : (counter_2  ? ((~counter_1  & (reg_2  ? ((~reg_4  & (((~reg_1  ^ reg_6 ) & (reg_3  ? (~reg_7  ^ reg_8 ) : (~reg_7  & ~reg_8 ))) | (~reg_1  & reg_7  & (reg_3  ? (reg_6  & reg_8 ) : (~reg_6  & ~reg_8 ))))) | (~reg_1  & reg_4  & ((~reg_3  & ~reg_6  & ~reg_7  & ~reg_8 ) | (reg_3  & (reg_6  ? (reg_7  & reg_8 ) : (~reg_7  & ~reg_8 )))))) : ((reg_4  & (reg_1  ? (~reg_3  & (reg_6  ? (~reg_7  & ~reg_8 ) : (reg_7  & reg_8 ))) : (reg_3  & (reg_6  ? reg_8  : (~reg_7  & ~reg_8 ))))) | (~reg_3  & ~reg_4  & reg_7  & reg_8  & (~reg_1  | (reg_1  & ~reg_6 )))))) | (~reg_2  & reg_3  & counter_1  & reg_1  & reg_7  & ~reg_8  & reg_4  & ~reg_6 )) : (reg_3  ? ((~reg_7  & ((~reg_8  & ((~reg_6  & ((counter_1  & ~reg_2  & reg_4 ) | (~counter_1  & reg_2  & ~reg_4 ) | (~counter_1  & ~reg_1  & ~reg_2  & ~reg_4 ))) | (reg_1  & ~reg_2  & reg_6  & (counter_1  ^ reg_4 )))) | (~counter_1  & reg_1  & ~reg_2  & ~reg_4  & ~reg_6  & reg_8 ))) | (~counter_1  & ~reg_4  & reg_7  & reg_8  & (reg_1  ? (~reg_2  ^ reg_6 ) : (reg_2  & reg_6 )))) : (reg_6  ? (counter_1  ? (reg_1  ? ((~reg_2  & ~reg_4  & reg_7  & reg_8 ) | (reg_2  & reg_4  & ~reg_7  & ~reg_8 )) : ((~reg_2  & reg_4  & reg_7  & reg_8 ) | (reg_2  & ~reg_4  & ~reg_7  & ~reg_8 ))) : ((~reg_4  & ((reg_7  & (reg_1  ? (~reg_2  ^ reg_8 ) : (~reg_2  & reg_8 ))) | (~reg_1  & ~reg_7  & (reg_2  ^ reg_8 )))) | (~reg_1  & reg_2  & reg_4  & reg_7  & ~reg_8 ))) : ((reg_2  & ((reg_1  & ((counter_1  & ~reg_4  & (~reg_7  ^ reg_8 )) | (reg_7  & reg_8  & ~counter_1  & reg_4 ))) | (~counter_1  & ~reg_1  & ~reg_4  & ~reg_7  & ~reg_8 ))) | (~counter_1  & ~reg_1  & ~reg_2  & ~reg_4  & ~reg_7  & reg_8 )))))) : (reg_0  ? (reg_1  ? ((~counter_2  & ~reg_7  & ~reg_8  & ((counter_1  & ~reg_3  & (reg_4  ^ reg_6 )) | (~reg_4  & reg_6  & ~counter_1  & reg_3 ))) | (~counter_1  & counter_2  & reg_7  & reg_8  & (reg_3  ? (~reg_4  & reg_6 ) : (reg_4  & ~reg_6 ))) | (reg_7  & ((~reg_4  & ((~counter_2  & ((reg_8  & ((counter_1  & (reg_2  ? (~reg_3  & ~reg_6 ) : (reg_3  & reg_6 ))) | (~counter_1  & reg_2  & reg_3  & reg_6 ))) | (~counter_1  & reg_2  & reg_3  & ~reg_6  & ~reg_8 ))) | (~counter_1  & counter_2  & ((~reg_2  & (reg_3  ? (~reg_6  & ~reg_8 ) : (reg_6  & reg_8 ))) | (reg_2  & ~reg_3  & reg_6  & ~reg_8 ))))) | (~counter_1  & reg_4  & ((counter_2  & ((reg_2  & reg_8  & (reg_3  ^ reg_6 )) | (~reg_2  & reg_3  & reg_6  & ~reg_8 ))) | (~counter_2  & ~reg_2  & reg_3  & ~reg_6  & reg_8 ))))) | (~counter_1  & ~reg_7  & ~reg_8  & ((counter_2  & ((~reg_2  & ~reg_4  & (~reg_3  ^ reg_6 )) | (reg_2  & reg_3  & reg_4  & ~reg_6 ))) | (~counter_2  & ~reg_2  & ~reg_3  & reg_4  & ~reg_6 )))) : (((reg_2  ? (reg_3  & reg_6 ) : (~reg_3  & ~reg_6 )) & ((counter_1  & ~counter_2  & ~reg_4  & reg_7  & reg_8 ) | (~counter_1  & counter_2  & reg_4  & ~reg_7  & ~reg_8 ))) | (~counter_1  & (reg_2  ? ((reg_6  & (((reg_3  ^ reg_4 ) & (counter_2  ? (reg_7  & reg_8 ) : (~reg_7  & ~reg_8 ))) | (~counter_2  & reg_3  & reg_4  & reg_7  & reg_8 ))) | (~counter_2  & ~reg_6  & ((reg_3  & (reg_4  ? (~reg_7  & reg_8 ) : (reg_7  & ~reg_8 ))) | (~reg_3  & reg_4  & ~reg_7  & ~reg_8 )))) : ((~reg_4  & (counter_2  ? (reg_3  & (reg_6  ? (~reg_7  & ~reg_8 ) : (reg_7  & reg_8 ))) : (~reg_3  & reg_8  & (reg_6  ^ reg_7 )))) | (~counter_2  & ~reg_3  & reg_4  & ~reg_6  & reg_7  & ~reg_8 )))))) : ((~counter_1  & reg_7  & reg_8  & ((~reg_1  & reg_2  & (counter_2  ? reg_6  : (~reg_3  & ~reg_6 ))) | (~counter_2  & reg_1  & ~reg_2  & ~reg_3  & reg_6 ))) | (~reg_1  & reg_2  & counter_1  & ~counter_2  & reg_3  & reg_6  & ~reg_7  & ~reg_8 ) | (reg_8  & ((reg_7  & ((~reg_3  & ((reg_1  & ((reg_4  & ((~reg_6  & (counter_1  ? (counter_2  ^ reg_2 ) : (counter_2  & reg_2 ))) | (~counter_1  & ~counter_2  & reg_2  & reg_6 ))) | (~counter_1  & ~counter_2  & reg_2  & ~reg_4  & ~reg_6 ))) | (~counter_1  & ~counter_2  & ~reg_1  & (reg_2  ? (~reg_4  & reg_6 ) : (~reg_4  ^ reg_6 ))))) | (~counter_1  & ~reg_2  & reg_3  & ~reg_4  & ((reg_1  & ~reg_6 ) | (~reg_1  & reg_6 ) | (counter_2  & ~reg_1  & ~reg_6 ))))) | (~counter_1  & ~reg_7  & ((reg_3  & ((~reg_1  & ((reg_6  & (counter_2  ? (~reg_2  ^ reg_4 ) : (~reg_2  & reg_4 ))) | (~counter_2  & reg_2  & ~reg_4  & ~reg_6 ))) | (~counter_2  & reg_1  & reg_2  & ~reg_4  & reg_6 ))) | (~reg_3  & reg_4  & reg_6  & ~counter_2  & reg_1  & reg_2 ))))) | (~reg_8  & ((~reg_7  & ((reg_1  & ((~counter_2  & ~reg_2  & ((counter_1  & (reg_3  ? (~reg_4  & ~reg_6 ) : (reg_4  & reg_6 ))) | (reg_4  & ~reg_6  & ~counter_1  & ~reg_3 ))) | (~counter_1  & counter_2  & reg_2  & reg_3  & (reg_4  ^ reg_6 )))) | (~counter_1  & ~reg_1  & ((reg_2  & ((counter_2  & ~reg_6  & (reg_3  ^ reg_4 )) | (~counter_2  & reg_3  & reg_4  & reg_6 ))) | (counter_2  & ~reg_2  & ~reg_3  & reg_4  & ~reg_6 ))))) | (~reg_1  & ~reg_2  & ~counter_1  & ~counter_2  & reg_6  & reg_7  & ~reg_3  & ~reg_4 )))))) : ((((reg_5  & reg_7  & reg_8  & reg_3  & reg_4 ) | (~reg_5  & ~reg_7  & ~reg_8  & ~reg_3  & ~reg_4 )) & ((~reg_1  & reg_6  & ((counter_1  & ~counter_2  & (reg_0  ^ reg_2 )) | (~counter_1  & counter_2  & reg_0  & reg_2 ))) | (~counter_1  & counter_2  & reg_0  & reg_1  & ~reg_2  & ~reg_6 ))) | (counter_2  & (reg_0  ? (reg_1  ? ((reg_5  & ((reg_7  & (counter_1  ? ((~reg_2  & reg_3  & ~reg_4  & ~reg_6  & reg_8 ) | (reg_2  & ~reg_3  & reg_4  & reg_6  & ~reg_8 )) : (~reg_2  & ((reg_3  & reg_6  & (reg_4  ^ ~reg_8 )) | (~reg_6  & reg_8  & ~reg_3  & ~reg_4 ))))) | (~counter_1  & ~reg_7  & ((reg_2  & ~reg_3  & reg_4  & reg_6  & ~reg_8 ) | (~reg_2  & ~reg_4  & ~reg_6  & (~reg_3  ^ ~reg_8 )))))) | (~counter_1  & ~reg_5  & ~reg_6  & ((reg_3  & ((~reg_2  & reg_4  & reg_7  & reg_8 ) | (reg_2  & ~reg_4  & ~reg_7  & ~reg_8 ))) | (reg_2  & ~reg_3  & ~reg_7  & ~reg_8 )))) : ((reg_5  & ((~reg_2  & ((~counter_1  & ~reg_4  & ~reg_6  & ~reg_8  & (~reg_3  ^ reg_7 )) | (reg_6  & reg_7  & reg_8  & counter_1  & reg_3  & reg_4 ))) | (reg_4  & ~reg_6  & ~reg_7  & ~reg_8  & ~counter_1  & reg_2  & ~reg_3 ))) | (~reg_4  & ~reg_5  & ((~reg_6  & (counter_1  ? ((~reg_2  & reg_3  & reg_7  & reg_8 ) | (reg_2  & ~reg_3  & ~reg_7  & ~reg_8 )) : ((reg_2  & reg_7  & reg_8 ) | (~reg_2  & ~reg_3  & ~reg_7  & ~reg_8 )))) | (reg_6  & ~reg_7  & ~reg_8  & counter_1  & reg_2  & reg_3 ))))) : ((reg_4  & ((~reg_6  & (((reg_2  ? (~reg_7  & ~reg_8 ) : (reg_7  & reg_8 )) & ((reg_3  & reg_5  & counter_1  & reg_1 ) | (~counter_1  & ~reg_1  & ~reg_3  & ~reg_5 ))) | (~counter_1  & (reg_1  ? (reg_2  ? ((~reg_3  & (reg_5  ? (reg_7  & reg_8 ) : (~reg_7  & ~reg_8 ))) | (reg_3  & ~reg_5  & ~reg_7  & ~reg_8 )) : ((~reg_7  & reg_8  & ~reg_3  & ~reg_5 ) | (reg_7  & ~reg_8  & reg_3  & reg_5 ))) : (~reg_3  & ((~reg_2  & ~reg_7  & (reg_5  ^ ~reg_8 )) | (reg_2  & reg_5  & reg_7  & reg_8 ))))) | (counter_1  & ~reg_1  & reg_2  & ~reg_3  & ~reg_5  & ~reg_7  & ~reg_8 ))) | (~counter_1  & reg_6  & (reg_3  ? (reg_5  & ((~reg_1  & reg_2  & (~reg_7  ^ reg_8 )) | (reg_1  & ~reg_2  & ~reg_7  & ~reg_8 ))) : ((~reg_2  & ((~reg_1  & ~reg_5  & ~reg_7  & ~reg_8 ) | (reg_1  & (reg_5  ? (reg_7  & reg_8 ) : (~reg_7  & ~reg_8 ))))) | (~reg_1  & reg_2  & (reg_5  ? (~reg_7  & ~reg_8 ) : (reg_7  & reg_8 )))))))) | (~counter_1  & ~reg_4  & (reg_2  ? ((reg_6  & ((reg_1  & ~reg_8  & (reg_3  ? (~reg_5  & reg_7 ) : (reg_5  & ~reg_7 ))) | (~reg_1  & reg_3  & reg_5  & reg_7  & reg_8 ))) | (~reg_1  & ~reg_6  & reg_8  & (reg_3  ? (reg_5  & reg_7 ) : ~reg_7 ))) : ((reg_6  & ((~reg_1  & ~reg_5  & reg_7  & reg_8 ) | (reg_1  & reg_5  & ~reg_7  & ~reg_8 ) | (~reg_1  & reg_3  & reg_5  & ~reg_7  & ~reg_8 ))) | (reg_5  & ~reg_6  & ((~reg_1  & (reg_3  ? (reg_7  & reg_8 ) : (~reg_7  & ~reg_8 ))) | (reg_1  & ~reg_3  & ~reg_7  & ~reg_8 ))))))))) | (counter_1  & ~counter_2  & (reg_7  ? (reg_5  ? (reg_1  ? ((reg_8  & (reg_0  ? (reg_6  & (reg_2  ? (~reg_3  & reg_4 ) : (reg_3  & ~reg_4 ))) : (reg_3  & ~reg_6  & (~reg_2  | (reg_2  & ~reg_4 ))))) | (~reg_0  & reg_2  & ~reg_3  & ~reg_8  & (reg_4  ^ reg_6 ))) : (reg_4  & reg_8  & ((reg_0  & (reg_2  ? (reg_3  & ~reg_6 ) : (~reg_3  & reg_6 ))) | (~reg_0  & reg_2  & ~reg_3  & ~reg_6 )))) : (reg_0  ? (reg_2  ? (~reg_6  & reg_8  & (~reg_1  ^ ~reg_4 )) : ((reg_1  & (reg_3  ? (reg_4  ? (reg_6  & ~reg_8 ) : (~reg_6  & reg_8 )) : (reg_6  & reg_8 ))) | (~reg_1  & ~reg_3  & reg_4  & ~reg_6  & ~reg_8 ))) : (reg_8  & ((~reg_2  & reg_3  & ~reg_4  & reg_6 ) | (reg_2  & ~reg_3  & reg_4  & ~reg_6 ) | (~reg_4  & ((reg_2  & (reg_1  ? ~reg_3  : (reg_3  & reg_6 ))) | (~reg_1  & ~reg_2  & reg_3  & ~reg_6 ))))))) : (reg_6  ? (reg_0  ? (~reg_8  & ((reg_4  & ((~reg_1  & reg_2  & (reg_3  | (~reg_3  & ~reg_5 ))) | (reg_1  & ~reg_2  & ~reg_3  & reg_5 ))) | (reg_2  & ~reg_4  & ~reg_5  & (reg_1  | (~reg_1  & reg_3 ))))) : ((reg_4  & ((reg_1  & ((~reg_2  & reg_3  & ~reg_5  & reg_8 ) | (reg_2  & ~reg_3  & reg_5  & ~reg_8 ))) | (~reg_1  & reg_2  & ~reg_3  & reg_5  & ~reg_8 ))) | (~reg_1  & ~reg_4  & ((~reg_2  & ~reg_3  & reg_5  & reg_8 ) | (reg_2  & reg_3  & ~reg_5  & ~reg_8 ))))) : (~reg_8  & ((reg_5  & ((~reg_0  & ~reg_1  & reg_2  & reg_3 ) | (reg_0  & reg_1  & ~reg_2  & ~reg_3 ) | (~reg_1  & ((reg_0  & (reg_2  ? (reg_3  & reg_4 ) : (~reg_3  & ~reg_4 ))) | (~reg_0  & ~reg_2  & reg_3  & ~reg_4 ))) | (~reg_0  & reg_1  & (reg_2  ? (reg_3  & ~reg_4 ) : (~reg_3  & reg_4 ))))) | (reg_0  & ~reg_1  & reg_2  & reg_3  & reg_4  & ~reg_5 ))))))))));
  assign out = n54_1 ? n96 : n97;
  always @ (posedge clock) begin
    reg_0  <= n24;
    reg_1  <= n29;
    reg_2  <= n34;
    reg_3  <= n39;
    reg_4  <= n44;
    reg_5  <= n49;
    reg_6  <= n54;
    reg_7  <= n59;
    reg_8  <= n64;
    counter_0  <= n69;
    counter_1  <= n74;
    counter_2  <= n79;
    counter_3  <= n84;
    counter_4  <= n89;
  end
  initial begin
    reg_0  <= 1'b0;
    reg_1  <= 1'b0;
    reg_2  <= 1'b0;
    reg_3  <= 1'b0;
    reg_4  <= 1'b0;
    reg_5  <= 1'b0;
    reg_6  <= 1'b0;
    reg_7  <= 1'b0;
    reg_8  <= 1'b0;
    counter_0  <= 1'b0;
    counter_1  <= 1'b0;
    counter_2  <= 1'b0;
    counter_3  <= 1'b0;
    counter_4  <= 1'b0;
  end
endmodule


