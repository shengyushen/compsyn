
module scrambler ( CLK, reset, data_66b_tpg, data_scrambled, 
        assertion_shengyushen );
  input [63:0] data_66b_tpg;
  output [63:0] data_scrambled;
  input CLK, reset;
  output assertion_shengyushen;
  wire   U4_Z_0, U4_Z_1, U4_Z_2, U4_Z_3, U4_Z_4, U4_Z_5, U4_Z_6, U4_Z_7,
         U4_Z_8, U4_Z_9, U4_Z_10, U4_Z_11, U4_Z_12, U4_Z_13, U4_Z_14, U4_Z_15,
         U4_Z_16, U4_Z_17, U4_Z_18, U4_Z_19, U4_Z_20, U4_Z_21, U4_Z_22,
         U4_Z_23, U4_Z_24, U4_Z_25, U4_Z_26, U4_Z_27, U4_Z_28, U4_Z_29,
         U4_Z_30, U4_Z_31, U4_Z_32, U4_Z_33, U4_Z_34, U4_Z_35, U4_Z_36,
         U4_Z_37, U4_Z_38, U4_Z_39, U4_Z_40, U4_Z_41, U4_Z_42, U4_Z_43,
         U4_Z_44, U4_Z_45, U4_Z_46, U4_Z_47, U4_Z_48, U4_Z_49, U4_Z_50,
         U4_Z_51, U4_Z_52, U4_Z_53, U4_Z_54, U4_Z_55, U4_Z_56, U4_Z_57, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303;
  wire   [181:124] n;

  IV I_0 ( .A(reset), .Z(assertion_shengyushen) );
  FD1 data_prev_reg_0_ ( .D(U4_Z_0), .CP(CLK), .Q(n[124]) );
  FD1 data_prev_reg_52_ ( .D(U4_Z_52), .CP(CLK), .Q(n[176]) );
  FD1 data_prev_reg_46_ ( .D(U4_Z_46), .CP(CLK), .Q(n[170]) );
  FD1 data_prev_reg_40_ ( .D(U4_Z_40), .CP(CLK), .Q(n[164]) );
  FD1 data_prev_reg_34_ ( .D(U4_Z_34), .CP(CLK), .Q(n[158]) );
  FD1 data_prev_reg_9_ ( .D(U4_Z_9), .CP(CLK), .Q(n[133]) );
  FD1 data_prev_reg_3_ ( .D(U4_Z_3), .CP(CLK), .Q(n[127]) );
  FD1 data_prev_reg_55_ ( .D(U4_Z_55), .CP(CLK), .Q(n[179]) );
  FD1 data_prev_reg_49_ ( .D(U4_Z_49), .CP(CLK), .Q(n[173]) );
  FD1 data_prev_reg_43_ ( .D(U4_Z_43), .CP(CLK), .Q(n[167]) );
  FD1 data_prev_reg_37_ ( .D(U4_Z_37), .CP(CLK), .Q(n[161]) );
  FD1 data_prev_reg_31_ ( .D(U4_Z_31), .CP(CLK), .Q(n[155]) );
  FD1 data_prev_reg_6_ ( .D(U4_Z_6), .CP(CLK), .Q(n[130]) );
  FD1 data_prev_reg_39_ ( .D(U4_Z_39), .CP(CLK), .Q(n[163]) );
  FD1 data_prev_reg_33_ ( .D(U4_Z_33), .CP(CLK), .Q(n[157]) );
  FD1 data_prev_reg_27_ ( .D(U4_Z_27), .CP(CLK), .Q(n[151]) );
  FD1 data_prev_reg_21_ ( .D(U4_Z_21), .CP(CLK), .Q(n[145]) );
  FD1 data_prev_reg_15_ ( .D(U4_Z_15), .CP(CLK), .Q(n[139]) );
  FD1 data_prev_reg_8_ ( .D(U4_Z_8), .CP(CLK), .Q(n[132]) );
  FD1 data_prev_reg_2_ ( .D(U4_Z_2), .CP(CLK), .Q(n[126]) );
  FD1 data_prev_reg_54_ ( .D(U4_Z_54), .CP(CLK), .Q(n[178]) );
  FD1 data_prev_reg_48_ ( .D(U4_Z_48), .CP(CLK), .Q(n[172]) );
  FD1 data_prev_reg_42_ ( .D(U4_Z_42), .CP(CLK), .Q(n[166]) );
  FD1 data_prev_reg_36_ ( .D(U4_Z_36), .CP(CLK), .Q(n[160]) );
  FD1 data_prev_reg_30_ ( .D(U4_Z_30), .CP(CLK), .Q(n[154]) );
  FD1 data_prev_reg_24_ ( .D(U4_Z_24), .CP(CLK), .Q(n[148]) );
  FD1 data_prev_reg_18_ ( .D(U4_Z_18), .CP(CLK), .Q(n[142]) );
  FD1 data_prev_reg_12_ ( .D(U4_Z_12), .CP(CLK), .Q(n[136]) );
  FD1 data_prev_reg_5_ ( .D(U4_Z_5), .CP(CLK), .Q(n[129]) );
  FD1 data_prev_reg_57_ ( .D(U4_Z_57), .CP(CLK), .Q(n[181]) );
  FD1 data_prev_reg_51_ ( .D(U4_Z_51), .CP(CLK), .Q(n[175]) );
  FD1 data_prev_reg_45_ ( .D(U4_Z_45), .CP(CLK), .Q(n[169]) );
  FD1 data_prev_reg_20_ ( .D(U4_Z_20), .CP(CLK), .Q(n[144]) );
  FD1 data_prev_reg_14_ ( .D(U4_Z_14), .CP(CLK), .Q(n[138]) );
  FD1 data_prev_reg_53_ ( .D(U4_Z_53), .CP(CLK), .Q(n[177]) );
  FD1 data_prev_reg_28_ ( .D(U4_Z_28), .CP(CLK), .Q(n[152]) );
  FD1 data_prev_reg_47_ ( .D(U4_Z_47), .CP(CLK), .Q(n[171]) );
  FD1 data_prev_reg_22_ ( .D(U4_Z_22), .CP(CLK), .Q(n[146]) );
  FD1 data_prev_reg_41_ ( .D(U4_Z_41), .CP(CLK), .Q(n[165]) );
  FD1 data_prev_reg_16_ ( .D(U4_Z_16), .CP(CLK), .Q(n[140]) );
  FD1 data_prev_reg_35_ ( .D(U4_Z_35), .CP(CLK), .Q(n[159]) );
  FD1 data_prev_reg_10_ ( .D(U4_Z_10), .CP(CLK), .Q(n[134]) );
  FD1 data_prev_reg_29_ ( .D(U4_Z_29), .CP(CLK), .Q(n[153]) );
  FD1 data_prev_reg_23_ ( .D(U4_Z_23), .CP(CLK), .Q(n[147]) );
  FD1 data_prev_reg_17_ ( .D(U4_Z_17), .CP(CLK), .Q(n[141]) );
  FD1 data_prev_reg_11_ ( .D(U4_Z_11), .CP(CLK), .Q(n[135]) );
  FD1 data_prev_reg_4_ ( .D(U4_Z_4), .CP(CLK), .Q(n[128]) );
  FD1 data_prev_reg_56_ ( .D(U4_Z_56), .CP(CLK), .Q(n[180]) );
  FD1 data_prev_reg_50_ ( .D(U4_Z_50), .CP(CLK), .Q(n[174]) );
  FD1 data_prev_reg_25_ ( .D(U4_Z_25), .CP(CLK), .Q(n[149]) );
  FD1 data_prev_reg_44_ ( .D(U4_Z_44), .CP(CLK), .Q(n[168]) );
  FD1 data_prev_reg_19_ ( .D(U4_Z_19), .CP(CLK), .Q(n[143]) );
  FD1 data_prev_reg_38_ ( .D(U4_Z_38), .CP(CLK), .Q(n[162]) );
  FD1 data_prev_reg_13_ ( .D(U4_Z_13), .CP(CLK), .Q(n[137]) );
  FD1 data_prev_reg_32_ ( .D(U4_Z_32), .CP(CLK), .Q(n[156]) );
  FD1 data_prev_reg_26_ ( .D(U4_Z_26), .CP(CLK), .Q(n[150]) );
  FD1 data_prev_reg_7_ ( .D(U4_Z_7), .CP(CLK), .Q(n[131]) );
  FD1 data_prev_reg_1_ ( .D(U4_Z_1), .CP(CLK), .Q(n[125]) );
  IV U164 ( .A(data_66b_tpg[63]), .Z(n477) );
  IV U165 ( .A(data_66b_tpg[62]), .Z(n478) );
  IV U166 ( .A(data_66b_tpg[61]), .Z(n479) );
  IV U167 ( .A(data_66b_tpg[60]), .Z(n480) );
  IV U168 ( .A(data_66b_tpg[59]), .Z(n481) );
  IV U169 ( .A(data_66b_tpg[58]), .Z(n482) );
  IV U170 ( .A(data_66b_tpg[24]), .Z(n483) );
  IV U171 ( .A(data_66b_tpg[23]), .Z(n484) );
  IV U172 ( .A(data_66b_tpg[22]), .Z(n485) );
  IV U173 ( .A(data_66b_tpg[21]), .Z(n486) );
  IV U174 ( .A(data_66b_tpg[20]), .Z(n487) );
  IV U175 ( .A(data_66b_tpg[19]), .Z(n488) );
  AN2 U618 ( .A(assertion_shengyushen), .B(data_scrambled[15]), .Z(U4_Z_9) );
  AN2 U619 ( .A(assertion_shengyushen), .B(data_scrambled[14]), .Z(U4_Z_8) );
  AN2 U620 ( .A(assertion_shengyushen), .B(data_scrambled[13]), .Z(U4_Z_7) );
  AN2 U621 ( .A(assertion_shengyushen), .B(data_scrambled[12]), .Z(U4_Z_6) );
  AN2 U622 ( .A(assertion_shengyushen), .B(data_scrambled[63]), .Z(U4_Z_57) );
  AN2 U623 ( .A(assertion_shengyushen), .B(data_scrambled[62]), .Z(U4_Z_56) );
  AN2 U624 ( .A(assertion_shengyushen), .B(data_scrambled[61]), .Z(U4_Z_55) );
  AN2 U625 ( .A(assertion_shengyushen), .B(data_scrambled[60]), .Z(U4_Z_54) );
  AN2 U626 ( .A(assertion_shengyushen), .B(data_scrambled[59]), .Z(U4_Z_53) );
  AN2 U627 ( .A(assertion_shengyushen), .B(data_scrambled[58]), .Z(U4_Z_52) );
  AN2 U628 ( .A(assertion_shengyushen), .B(data_scrambled[57]), .Z(U4_Z_51) );
  AN2 U629 ( .A(assertion_shengyushen), .B(data_scrambled[56]), .Z(U4_Z_50) );
  AN2 U630 ( .A(assertion_shengyushen), .B(data_scrambled[11]), .Z(U4_Z_5) );
  AN2 U631 ( .A(assertion_shengyushen), .B(data_scrambled[55]), .Z(U4_Z_49) );
  AN2 U632 ( .A(assertion_shengyushen), .B(data_scrambled[54]), .Z(U4_Z_48) );
  AN2 U633 ( .A(assertion_shengyushen), .B(data_scrambled[53]), .Z(U4_Z_47) );
  AN2 U634 ( .A(assertion_shengyushen), .B(data_scrambled[52]), .Z(U4_Z_46) );
  AN2 U635 ( .A(assertion_shengyushen), .B(data_scrambled[51]), .Z(U4_Z_45) );
  AN2 U636 ( .A(assertion_shengyushen), .B(data_scrambled[50]), .Z(U4_Z_44) );
  AN2 U637 ( .A(assertion_shengyushen), .B(data_scrambled[49]), .Z(U4_Z_43) );
  AN2 U638 ( .A(assertion_shengyushen), .B(data_scrambled[48]), .Z(U4_Z_42) );
  AN2 U639 ( .A(assertion_shengyushen), .B(data_scrambled[47]), .Z(U4_Z_41) );
  AN2 U640 ( .A(assertion_shengyushen), .B(data_scrambled[46]), .Z(U4_Z_40) );
  AN2 U641 ( .A(assertion_shengyushen), .B(data_scrambled[10]), .Z(U4_Z_4) );
  AN2 U642 ( .A(assertion_shengyushen), .B(data_scrambled[45]), .Z(U4_Z_39) );
  AN2 U643 ( .A(assertion_shengyushen), .B(data_scrambled[44]), .Z(U4_Z_38) );
  AN2 U644 ( .A(assertion_shengyushen), .B(data_scrambled[43]), .Z(U4_Z_37) );
  AN2 U645 ( .A(assertion_shengyushen), .B(data_scrambled[42]), .Z(U4_Z_36) );
  AN2 U646 ( .A(assertion_shengyushen), .B(data_scrambled[41]), .Z(U4_Z_35) );
  AN2 U647 ( .A(assertion_shengyushen), .B(data_scrambled[40]), .Z(U4_Z_34) );
  AN2 U648 ( .A(assertion_shengyushen), .B(data_scrambled[39]), .Z(U4_Z_33) );
  AN2 U649 ( .A(assertion_shengyushen), .B(data_scrambled[38]), .Z(U4_Z_32) );
  AN2 U650 ( .A(assertion_shengyushen), .B(data_scrambled[37]), .Z(U4_Z_31) );
  AN2 U651 ( .A(assertion_shengyushen), .B(data_scrambled[36]), .Z(U4_Z_30) );
  AN2 U652 ( .A(assertion_shengyushen), .B(data_scrambled[9]), .Z(U4_Z_3) );
  AN2 U653 ( .A(assertion_shengyushen), .B(data_scrambled[35]), .Z(U4_Z_29) );
  AN2 U654 ( .A(assertion_shengyushen), .B(data_scrambled[34]), .Z(U4_Z_28) );
  AN2 U655 ( .A(assertion_shengyushen), .B(data_scrambled[33]), .Z(U4_Z_27) );
  AN2 U656 ( .A(assertion_shengyushen), .B(data_scrambled[32]), .Z(U4_Z_26) );
  AN2 U657 ( .A(assertion_shengyushen), .B(data_scrambled[31]), .Z(U4_Z_25) );
  AN2 U658 ( .A(assertion_shengyushen), .B(data_scrambled[30]), .Z(U4_Z_24) );
  AN2 U659 ( .A(assertion_shengyushen), .B(data_scrambled[29]), .Z(U4_Z_23) );
  AN2 U660 ( .A(assertion_shengyushen), .B(data_scrambled[28]), .Z(U4_Z_22) );
  AN2 U661 ( .A(assertion_shengyushen), .B(data_scrambled[27]), .Z(U4_Z_21) );
  AN2 U662 ( .A(assertion_shengyushen), .B(data_scrambled[26]), .Z(U4_Z_20) );
  AN2 U663 ( .A(assertion_shengyushen), .B(data_scrambled[8]), .Z(U4_Z_2) );
  AN2 U664 ( .A(assertion_shengyushen), .B(data_scrambled[25]), .Z(U4_Z_19) );
  AN2 U665 ( .A(data_scrambled[24]), .B(assertion_shengyushen), .Z(U4_Z_18) );
  AN2 U666 ( .A(data_scrambled[23]), .B(assertion_shengyushen), .Z(U4_Z_17) );
  AN2 U667 ( .A(data_scrambled[22]), .B(assertion_shengyushen), .Z(U4_Z_16) );
  AN2 U668 ( .A(data_scrambled[21]), .B(assertion_shengyushen), .Z(U4_Z_15) );
  AN2 U669 ( .A(data_scrambled[20]), .B(assertion_shengyushen), .Z(U4_Z_14) );
  AN2 U670 ( .A(data_scrambled[19]), .B(assertion_shengyushen), .Z(U4_Z_13) );
  AN2 U671 ( .A(assertion_shengyushen), .B(data_scrambled[18]), .Z(U4_Z_12) );
  AN2 U672 ( .A(assertion_shengyushen), .B(data_scrambled[17]), .Z(U4_Z_11) );
  AN2 U673 ( .A(assertion_shengyushen), .B(data_scrambled[16]), .Z(U4_Z_10) );
  AN2 U674 ( .A(assertion_shengyushen), .B(data_scrambled[7]), .Z(U4_Z_1) );
  AN2 U675 ( .A(assertion_shengyushen), .B(data_scrambled[6]), .Z(U4_Z_0) );
  OR2 U676 ( .A(n811), .B(n812), .Z(data_scrambled[63]) );
  AN2 U677 ( .A(n813), .B(data_scrambled[24]), .Z(n812) );
  IV U678 ( .A(n814), .Z(n811) );
  OR2 U679 ( .A(data_scrambled[24]), .B(n813), .Z(n814) );
  OR2 U680 ( .A(n815), .B(n816), .Z(n813) );
  AN2 U681 ( .A(data_scrambled[5]), .B(n817), .Z(n816) );
  IV U682 ( .A(n477), .Z(n817) );
  AN2 U683 ( .A(n477), .B(n818), .Z(n815) );
  OR2 U684 ( .A(n819), .B(n820), .Z(data_scrambled[62]) );
  AN2 U685 ( .A(n821), .B(data_scrambled[23]), .Z(n820) );
  IV U686 ( .A(n822), .Z(n819) );
  OR2 U687 ( .A(data_scrambled[23]), .B(n821), .Z(n822) );
  OR2 U688 ( .A(n823), .B(n824), .Z(n821) );
  AN2 U689 ( .A(data_scrambled[4]), .B(n825), .Z(n824) );
  IV U690 ( .A(n478), .Z(n825) );
  AN2 U691 ( .A(n478), .B(n826), .Z(n823) );
  OR2 U692 ( .A(n827), .B(n828), .Z(data_scrambled[61]) );
  AN2 U693 ( .A(n829), .B(data_scrambled[22]), .Z(n828) );
  IV U694 ( .A(n830), .Z(n827) );
  OR2 U695 ( .A(data_scrambled[22]), .B(n829), .Z(n830) );
  OR2 U696 ( .A(n831), .B(n832), .Z(n829) );
  AN2 U697 ( .A(data_scrambled[3]), .B(n833), .Z(n832) );
  IV U698 ( .A(n479), .Z(n833) );
  AN2 U699 ( .A(n479), .B(n834), .Z(n831) );
  OR2 U700 ( .A(n835), .B(n836), .Z(data_scrambled[60]) );
  AN2 U701 ( .A(n837), .B(data_scrambled[21]), .Z(n836) );
  IV U702 ( .A(n838), .Z(n835) );
  OR2 U703 ( .A(data_scrambled[21]), .B(n837), .Z(n838) );
  OR2 U704 ( .A(n839), .B(n840), .Z(n837) );
  AN2 U705 ( .A(data_scrambled[2]), .B(n841), .Z(n840) );
  IV U706 ( .A(n480), .Z(n841) );
  AN2 U707 ( .A(n480), .B(n842), .Z(n839) );
  OR2 U708 ( .A(n843), .B(n844), .Z(data_scrambled[59]) );
  AN2 U709 ( .A(n845), .B(data_scrambled[20]), .Z(n844) );
  IV U710 ( .A(n846), .Z(n843) );
  OR2 U711 ( .A(data_scrambled[20]), .B(n845), .Z(n846) );
  OR2 U712 ( .A(n847), .B(n848), .Z(n845) );
  AN2 U713 ( .A(data_scrambled[1]), .B(n849), .Z(n848) );
  IV U714 ( .A(n481), .Z(n849) );
  AN2 U715 ( .A(n481), .B(n850), .Z(n847) );
  OR2 U716 ( .A(n851), .B(n852), .Z(data_scrambled[58]) );
  AN2 U717 ( .A(n853), .B(data_scrambled[19]), .Z(n852) );
  IV U718 ( .A(n854), .Z(n851) );
  OR2 U719 ( .A(data_scrambled[19]), .B(n853), .Z(n854) );
  OR2 U720 ( .A(n855), .B(n856), .Z(n853) );
  AN2 U721 ( .A(data_scrambled[0]), .B(n857), .Z(n856) );
  IV U722 ( .A(n482), .Z(n857) );
  AN2 U723 ( .A(n482), .B(n858), .Z(n855) );
  OR2 U724 ( .A(n859), .B(n860), .Z(data_scrambled[57]) );
  IV U725 ( .A(n861), .Z(n860) );
  OR2 U726 ( .A(n862), .B(data_scrambled[18]), .Z(n861) );
  AN2 U727 ( .A(data_scrambled[18]), .B(n862), .Z(n859) );
  AN2 U728 ( .A(n863), .B(n864), .Z(n862) );
  OR2 U729 ( .A(n865), .B(n[181]), .Z(n864) );
  IV U730 ( .A(data_66b_tpg[57]), .Z(n865) );
  OR2 U731 ( .A(n866), .B(data_66b_tpg[57]), .Z(n863) );
  OR2 U732 ( .A(n867), .B(n868), .Z(data_scrambled[56]) );
  IV U733 ( .A(n869), .Z(n868) );
  OR2 U734 ( .A(n870), .B(data_scrambled[17]), .Z(n869) );
  AN2 U735 ( .A(data_scrambled[17]), .B(n870), .Z(n867) );
  AN2 U736 ( .A(n871), .B(n872), .Z(n870) );
  OR2 U737 ( .A(n873), .B(n[180]), .Z(n872) );
  IV U738 ( .A(data_66b_tpg[56]), .Z(n873) );
  OR2 U739 ( .A(n874), .B(data_66b_tpg[56]), .Z(n871) );
  OR2 U740 ( .A(n875), .B(n876), .Z(data_scrambled[55]) );
  IV U741 ( .A(n877), .Z(n876) );
  OR2 U742 ( .A(n878), .B(data_scrambled[16]), .Z(n877) );
  AN2 U743 ( .A(data_scrambled[16]), .B(n878), .Z(n875) );
  AN2 U744 ( .A(n879), .B(n880), .Z(n878) );
  OR2 U745 ( .A(n881), .B(n[179]), .Z(n880) );
  IV U746 ( .A(data_66b_tpg[55]), .Z(n881) );
  OR2 U747 ( .A(n882), .B(data_66b_tpg[55]), .Z(n879) );
  OR2 U748 ( .A(n883), .B(n884), .Z(data_scrambled[54]) );
  IV U749 ( .A(n885), .Z(n884) );
  OR2 U750 ( .A(n886), .B(data_scrambled[15]), .Z(n885) );
  AN2 U751 ( .A(data_scrambled[15]), .B(n886), .Z(n883) );
  AN2 U752 ( .A(n887), .B(n888), .Z(n886) );
  OR2 U753 ( .A(n889), .B(n[178]), .Z(n888) );
  IV U754 ( .A(data_66b_tpg[54]), .Z(n889) );
  OR2 U755 ( .A(n890), .B(data_66b_tpg[54]), .Z(n887) );
  OR2 U756 ( .A(n891), .B(n892), .Z(data_scrambled[15]) );
  IV U757 ( .A(n893), .Z(n892) );
  OR2 U758 ( .A(n894), .B(data_66b_tpg[15]), .Z(n893) );
  AN2 U759 ( .A(data_66b_tpg[15]), .B(n894), .Z(n891) );
  AN2 U760 ( .A(n895), .B(n896), .Z(n894) );
  OR2 U761 ( .A(n897), .B(n[158]), .Z(n896) );
  IV U762 ( .A(n[139]), .Z(n897) );
  OR2 U763 ( .A(n898), .B(n[139]), .Z(n895) );
  OR2 U764 ( .A(n899), .B(n900), .Z(data_scrambled[53]) );
  IV U765 ( .A(n901), .Z(n900) );
  OR2 U766 ( .A(n902), .B(data_scrambled[14]), .Z(n901) );
  AN2 U767 ( .A(data_scrambled[14]), .B(n902), .Z(n899) );
  AN2 U768 ( .A(n903), .B(n904), .Z(n902) );
  OR2 U769 ( .A(n905), .B(n[177]), .Z(n904) );
  IV U770 ( .A(data_66b_tpg[53]), .Z(n905) );
  OR2 U771 ( .A(n906), .B(data_66b_tpg[53]), .Z(n903) );
  OR2 U772 ( .A(n907), .B(n908), .Z(data_scrambled[14]) );
  IV U773 ( .A(n909), .Z(n908) );
  OR2 U774 ( .A(n910), .B(data_66b_tpg[14]), .Z(n909) );
  AN2 U775 ( .A(data_66b_tpg[14]), .B(n910), .Z(n907) );
  AN2 U776 ( .A(n911), .B(n912), .Z(n910) );
  OR2 U777 ( .A(n913), .B(n[157]), .Z(n912) );
  IV U778 ( .A(n[138]), .Z(n913) );
  OR2 U779 ( .A(n914), .B(n[138]), .Z(n911) );
  OR2 U780 ( .A(n915), .B(n916), .Z(data_scrambled[52]) );
  IV U781 ( .A(n917), .Z(n916) );
  OR2 U782 ( .A(n918), .B(data_scrambled[13]), .Z(n917) );
  AN2 U783 ( .A(data_scrambled[13]), .B(n918), .Z(n915) );
  AN2 U784 ( .A(n919), .B(n920), .Z(n918) );
  OR2 U785 ( .A(n921), .B(n[176]), .Z(n920) );
  IV U786 ( .A(data_66b_tpg[52]), .Z(n921) );
  OR2 U787 ( .A(n922), .B(data_66b_tpg[52]), .Z(n919) );
  OR2 U788 ( .A(n923), .B(n924), .Z(data_scrambled[13]) );
  IV U789 ( .A(n925), .Z(n924) );
  OR2 U790 ( .A(n926), .B(data_66b_tpg[13]), .Z(n925) );
  AN2 U791 ( .A(data_66b_tpg[13]), .B(n926), .Z(n923) );
  AN2 U792 ( .A(n927), .B(n928), .Z(n926) );
  OR2 U793 ( .A(n929), .B(n[156]), .Z(n928) );
  IV U794 ( .A(n[137]), .Z(n929) );
  OR2 U795 ( .A(n930), .B(n[137]), .Z(n927) );
  OR2 U796 ( .A(n931), .B(n932), .Z(data_scrambled[51]) );
  IV U797 ( .A(n933), .Z(n932) );
  OR2 U798 ( .A(n934), .B(data_scrambled[12]), .Z(n933) );
  AN2 U799 ( .A(data_scrambled[12]), .B(n934), .Z(n931) );
  AN2 U800 ( .A(n935), .B(n936), .Z(n934) );
  OR2 U801 ( .A(n937), .B(n[175]), .Z(n936) );
  IV U802 ( .A(data_66b_tpg[51]), .Z(n937) );
  OR2 U803 ( .A(n938), .B(data_66b_tpg[51]), .Z(n935) );
  OR2 U804 ( .A(n939), .B(n940), .Z(data_scrambled[12]) );
  IV U805 ( .A(n941), .Z(n940) );
  OR2 U806 ( .A(n942), .B(data_66b_tpg[12]), .Z(n941) );
  AN2 U807 ( .A(data_66b_tpg[12]), .B(n942), .Z(n939) );
  AN2 U808 ( .A(n943), .B(n944), .Z(n942) );
  OR2 U809 ( .A(n945), .B(n[155]), .Z(n944) );
  IV U810 ( .A(n[136]), .Z(n945) );
  OR2 U811 ( .A(n946), .B(n[136]), .Z(n943) );
  OR2 U812 ( .A(n947), .B(n948), .Z(data_scrambled[50]) );
  IV U813 ( .A(n949), .Z(n948) );
  OR2 U814 ( .A(n950), .B(data_scrambled[11]), .Z(n949) );
  AN2 U815 ( .A(data_scrambled[11]), .B(n950), .Z(n947) );
  AN2 U816 ( .A(n951), .B(n952), .Z(n950) );
  OR2 U817 ( .A(n953), .B(n[174]), .Z(n952) );
  IV U818 ( .A(data_66b_tpg[50]), .Z(n953) );
  OR2 U819 ( .A(n954), .B(data_66b_tpg[50]), .Z(n951) );
  OR2 U820 ( .A(n955), .B(n956), .Z(data_scrambled[11]) );
  IV U821 ( .A(n957), .Z(n956) );
  OR2 U822 ( .A(n958), .B(data_66b_tpg[11]), .Z(n957) );
  AN2 U823 ( .A(data_66b_tpg[11]), .B(n958), .Z(n955) );
  AN2 U824 ( .A(n959), .B(n960), .Z(n958) );
  OR2 U825 ( .A(n961), .B(n[154]), .Z(n960) );
  IV U826 ( .A(n[135]), .Z(n961) );
  OR2 U827 ( .A(n962), .B(n[135]), .Z(n959) );
  OR2 U828 ( .A(n963), .B(n964), .Z(data_scrambled[49]) );
  IV U829 ( .A(n965), .Z(n964) );
  OR2 U830 ( .A(n966), .B(data_scrambled[10]), .Z(n965) );
  AN2 U831 ( .A(data_scrambled[10]), .B(n966), .Z(n963) );
  AN2 U832 ( .A(n967), .B(n968), .Z(n966) );
  OR2 U833 ( .A(n969), .B(n[173]), .Z(n968) );
  IV U834 ( .A(data_66b_tpg[49]), .Z(n969) );
  OR2 U835 ( .A(n970), .B(data_66b_tpg[49]), .Z(n967) );
  OR2 U836 ( .A(n971), .B(n972), .Z(data_scrambled[48]) );
  IV U837 ( .A(n973), .Z(n972) );
  OR2 U838 ( .A(n974), .B(data_scrambled[9]), .Z(n973) );
  AN2 U839 ( .A(data_scrambled[9]), .B(n974), .Z(n971) );
  AN2 U840 ( .A(n975), .B(n976), .Z(n974) );
  OR2 U841 ( .A(n977), .B(n[172]), .Z(n976) );
  IV U842 ( .A(data_66b_tpg[48]), .Z(n977) );
  OR2 U843 ( .A(n978), .B(data_66b_tpg[48]), .Z(n975) );
  OR2 U844 ( .A(n979), .B(n980), .Z(data_scrambled[47]) );
  IV U845 ( .A(n981), .Z(n980) );
  OR2 U846 ( .A(n982), .B(data_scrambled[8]), .Z(n981) );
  AN2 U847 ( .A(data_scrambled[8]), .B(n982), .Z(n979) );
  AN2 U848 ( .A(n983), .B(n984), .Z(n982) );
  OR2 U849 ( .A(n985), .B(n[171]), .Z(n984) );
  IV U850 ( .A(data_66b_tpg[47]), .Z(n985) );
  OR2 U851 ( .A(n986), .B(data_66b_tpg[47]), .Z(n983) );
  OR2 U852 ( .A(n987), .B(n988), .Z(data_scrambled[46]) );
  IV U853 ( .A(n989), .Z(n988) );
  OR2 U854 ( .A(n990), .B(data_scrambled[7]), .Z(n989) );
  AN2 U855 ( .A(data_scrambled[7]), .B(n990), .Z(n987) );
  AN2 U856 ( .A(n991), .B(n992), .Z(n990) );
  OR2 U857 ( .A(n993), .B(n[170]), .Z(n992) );
  IV U858 ( .A(data_66b_tpg[46]), .Z(n993) );
  OR2 U859 ( .A(n994), .B(data_66b_tpg[46]), .Z(n991) );
  OR2 U860 ( .A(n995), .B(n996), .Z(data_scrambled[10]) );
  IV U861 ( .A(n997), .Z(n996) );
  OR2 U862 ( .A(n998), .B(data_66b_tpg[10]), .Z(n997) );
  AN2 U863 ( .A(data_66b_tpg[10]), .B(n998), .Z(n995) );
  AN2 U864 ( .A(n999), .B(n1000), .Z(n998) );
  OR2 U865 ( .A(n1001), .B(n[153]), .Z(n1000) );
  IV U866 ( .A(n[134]), .Z(n1001) );
  OR2 U867 ( .A(n1002), .B(n[134]), .Z(n999) );
  OR2 U868 ( .A(n1003), .B(n1004), .Z(data_scrambled[45]) );
  IV U869 ( .A(n1005), .Z(n1004) );
  OR2 U870 ( .A(n1006), .B(data_scrambled[6]), .Z(n1005) );
  AN2 U871 ( .A(data_scrambled[6]), .B(n1006), .Z(n1003) );
  AN2 U872 ( .A(n1007), .B(n1008), .Z(n1006) );
  OR2 U873 ( .A(n1009), .B(n[169]), .Z(n1008) );
  IV U874 ( .A(data_66b_tpg[45]), .Z(n1009) );
  OR2 U875 ( .A(n1010), .B(data_66b_tpg[45]), .Z(n1007) );
  OR2 U876 ( .A(n1011), .B(n1012), .Z(data_scrambled[44]) );
  IV U877 ( .A(n1013), .Z(n1012) );
  OR2 U878 ( .A(n1014), .B(data_scrambled[5]), .Z(n1013) );
  AN2 U879 ( .A(data_scrambled[5]), .B(n1014), .Z(n1011) );
  AN2 U880 ( .A(n1015), .B(n1016), .Z(n1014) );
  OR2 U881 ( .A(n1017), .B(n[168]), .Z(n1016) );
  IV U882 ( .A(data_66b_tpg[44]), .Z(n1017) );
  OR2 U883 ( .A(n1018), .B(data_66b_tpg[44]), .Z(n1015) );
  IV U884 ( .A(n818), .Z(data_scrambled[5]) );
  AN2 U885 ( .A(n1019), .B(n1020), .Z(n818) );
  OR2 U886 ( .A(n1021), .B(data_66b_tpg[5]), .Z(n1020) );
  IV U887 ( .A(n1022), .Z(n1019) );
  AN2 U888 ( .A(data_66b_tpg[5]), .B(n1021), .Z(n1022) );
  AN2 U889 ( .A(n1023), .B(n1024), .Z(n1021) );
  OR2 U890 ( .A(n1025), .B(n[148]), .Z(n1024) );
  IV U891 ( .A(n[129]), .Z(n1025) );
  OR2 U892 ( .A(n1026), .B(n[129]), .Z(n1023) );
  OR2 U893 ( .A(n1027), .B(n1028), .Z(data_scrambled[43]) );
  IV U894 ( .A(n1029), .Z(n1028) );
  OR2 U895 ( .A(n1030), .B(data_scrambled[4]), .Z(n1029) );
  AN2 U896 ( .A(data_scrambled[4]), .B(n1030), .Z(n1027) );
  AN2 U897 ( .A(n1031), .B(n1032), .Z(n1030) );
  OR2 U898 ( .A(n1033), .B(n[167]), .Z(n1032) );
  IV U899 ( .A(data_66b_tpg[43]), .Z(n1033) );
  OR2 U900 ( .A(n1034), .B(data_66b_tpg[43]), .Z(n1031) );
  IV U901 ( .A(n826), .Z(data_scrambled[4]) );
  AN2 U902 ( .A(n1035), .B(n1036), .Z(n826) );
  OR2 U903 ( .A(n1037), .B(data_66b_tpg[4]), .Z(n1036) );
  IV U904 ( .A(n1038), .Z(n1035) );
  AN2 U905 ( .A(data_66b_tpg[4]), .B(n1037), .Z(n1038) );
  AN2 U906 ( .A(n1039), .B(n1040), .Z(n1037) );
  OR2 U907 ( .A(n1041), .B(n[147]), .Z(n1040) );
  IV U908 ( .A(n[128]), .Z(n1041) );
  OR2 U909 ( .A(n1042), .B(n[128]), .Z(n1039) );
  OR2 U910 ( .A(n1043), .B(n1044), .Z(data_scrambled[42]) );
  IV U911 ( .A(n1045), .Z(n1044) );
  OR2 U912 ( .A(n1046), .B(data_scrambled[3]), .Z(n1045) );
  AN2 U913 ( .A(data_scrambled[3]), .B(n1046), .Z(n1043) );
  AN2 U914 ( .A(n1047), .B(n1048), .Z(n1046) );
  OR2 U915 ( .A(n1049), .B(n[166]), .Z(n1048) );
  IV U916 ( .A(data_66b_tpg[42]), .Z(n1049) );
  OR2 U917 ( .A(n1050), .B(data_66b_tpg[42]), .Z(n1047) );
  IV U918 ( .A(n834), .Z(data_scrambled[3]) );
  AN2 U919 ( .A(n1051), .B(n1052), .Z(n834) );
  OR2 U920 ( .A(n1053), .B(data_66b_tpg[3]), .Z(n1052) );
  IV U921 ( .A(n1054), .Z(n1051) );
  AN2 U922 ( .A(data_66b_tpg[3]), .B(n1053), .Z(n1054) );
  AN2 U923 ( .A(n1055), .B(n1056), .Z(n1053) );
  OR2 U924 ( .A(n1057), .B(n[146]), .Z(n1056) );
  IV U925 ( .A(n[127]), .Z(n1057) );
  OR2 U926 ( .A(n1058), .B(n[127]), .Z(n1055) );
  OR2 U927 ( .A(n1059), .B(n1060), .Z(data_scrambled[41]) );
  IV U928 ( .A(n1061), .Z(n1060) );
  OR2 U929 ( .A(n1062), .B(data_scrambled[2]), .Z(n1061) );
  AN2 U930 ( .A(data_scrambled[2]), .B(n1062), .Z(n1059) );
  AN2 U931 ( .A(n1063), .B(n1064), .Z(n1062) );
  OR2 U932 ( .A(n1065), .B(n[165]), .Z(n1064) );
  IV U933 ( .A(data_66b_tpg[41]), .Z(n1065) );
  OR2 U934 ( .A(n1066), .B(data_66b_tpg[41]), .Z(n1063) );
  IV U935 ( .A(n842), .Z(data_scrambled[2]) );
  AN2 U936 ( .A(n1067), .B(n1068), .Z(n842) );
  OR2 U937 ( .A(n1069), .B(data_66b_tpg[2]), .Z(n1068) );
  IV U938 ( .A(n1070), .Z(n1067) );
  AN2 U939 ( .A(data_66b_tpg[2]), .B(n1069), .Z(n1070) );
  AN2 U940 ( .A(n1071), .B(n1072), .Z(n1069) );
  OR2 U941 ( .A(n1073), .B(n[145]), .Z(n1072) );
  IV U942 ( .A(n[126]), .Z(n1073) );
  OR2 U943 ( .A(n1074), .B(n[126]), .Z(n1071) );
  OR2 U944 ( .A(n1075), .B(n1076), .Z(data_scrambled[40]) );
  IV U945 ( .A(n1077), .Z(n1076) );
  OR2 U946 ( .A(n1078), .B(data_scrambled[1]), .Z(n1077) );
  AN2 U947 ( .A(data_scrambled[1]), .B(n1078), .Z(n1075) );
  AN2 U948 ( .A(n1079), .B(n1080), .Z(n1078) );
  OR2 U949 ( .A(n1081), .B(n[164]), .Z(n1080) );
  IV U950 ( .A(data_66b_tpg[40]), .Z(n1081) );
  OR2 U951 ( .A(n1082), .B(data_66b_tpg[40]), .Z(n1079) );
  IV U952 ( .A(n850), .Z(data_scrambled[1]) );
  AN2 U953 ( .A(n1083), .B(n1084), .Z(n850) );
  OR2 U954 ( .A(n1085), .B(data_66b_tpg[1]), .Z(n1084) );
  IV U955 ( .A(n1086), .Z(n1083) );
  AN2 U956 ( .A(data_66b_tpg[1]), .B(n1085), .Z(n1086) );
  AN2 U957 ( .A(n1087), .B(n1088), .Z(n1085) );
  OR2 U958 ( .A(n1089), .B(n[144]), .Z(n1088) );
  IV U959 ( .A(n[125]), .Z(n1089) );
  OR2 U960 ( .A(n1090), .B(n[125]), .Z(n1087) );
  OR2 U961 ( .A(n1091), .B(n1092), .Z(data_scrambled[39]) );
  IV U962 ( .A(n1093), .Z(n1092) );
  OR2 U963 ( .A(n1094), .B(data_scrambled[0]), .Z(n1093) );
  AN2 U964 ( .A(data_scrambled[0]), .B(n1094), .Z(n1091) );
  AN2 U965 ( .A(n1095), .B(n1096), .Z(n1094) );
  OR2 U966 ( .A(n1097), .B(n[163]), .Z(n1096) );
  IV U967 ( .A(data_66b_tpg[39]), .Z(n1097) );
  OR2 U968 ( .A(n1098), .B(data_66b_tpg[39]), .Z(n1095) );
  IV U969 ( .A(n858), .Z(data_scrambled[0]) );
  AN2 U970 ( .A(n1099), .B(n1100), .Z(n858) );
  OR2 U971 ( .A(n1101), .B(data_66b_tpg[0]), .Z(n1100) );
  IV U972 ( .A(n1102), .Z(n1099) );
  AN2 U973 ( .A(data_66b_tpg[0]), .B(n1101), .Z(n1102) );
  AN2 U974 ( .A(n1103), .B(n1104), .Z(n1101) );
  OR2 U975 ( .A(n1105), .B(n[143]), .Z(n1104) );
  IV U976 ( .A(n[124]), .Z(n1105) );
  OR2 U977 ( .A(n1106), .B(n[124]), .Z(n1103) );
  OR2 U978 ( .A(n1107), .B(n1108), .Z(data_scrambled[38]) );
  AN2 U979 ( .A(n1109), .B(n1110), .Z(n1108) );
  IV U980 ( .A(n1111), .Z(n1107) );
  OR2 U981 ( .A(n1110), .B(n1109), .Z(n1111) );
  OR2 U982 ( .A(n1112), .B(n1113), .Z(n1109) );
  AN2 U983 ( .A(n[162]), .B(n866), .Z(n1113) );
  IV U984 ( .A(n[181]), .Z(n866) );
  AN2 U985 ( .A(n[181]), .B(n1114), .Z(n1112) );
  IV U986 ( .A(data_66b_tpg[38]), .Z(n1110) );
  OR2 U987 ( .A(n1115), .B(n1116), .Z(data_scrambled[37]) );
  AN2 U988 ( .A(n1117), .B(n1118), .Z(n1116) );
  IV U989 ( .A(n1119), .Z(n1115) );
  OR2 U990 ( .A(n1118), .B(n1117), .Z(n1119) );
  OR2 U991 ( .A(n1120), .B(n1121), .Z(n1117) );
  AN2 U992 ( .A(n[161]), .B(n874), .Z(n1121) );
  IV U993 ( .A(n[180]), .Z(n874) );
  AN2 U994 ( .A(n[180]), .B(n1122), .Z(n1120) );
  IV U995 ( .A(data_66b_tpg[37]), .Z(n1118) );
  OR2 U996 ( .A(n1123), .B(n1124), .Z(data_scrambled[36]) );
  AN2 U997 ( .A(n1125), .B(n1126), .Z(n1124) );
  IV U998 ( .A(n1127), .Z(n1123) );
  OR2 U999 ( .A(n1126), .B(n1125), .Z(n1127) );
  OR2 U1000 ( .A(n1128), .B(n1129), .Z(n1125) );
  AN2 U1001 ( .A(n[160]), .B(n882), .Z(n1129) );
  IV U1002 ( .A(n[179]), .Z(n882) );
  AN2 U1003 ( .A(n[179]), .B(n1130), .Z(n1128) );
  IV U1004 ( .A(data_66b_tpg[36]), .Z(n1126) );
  OR2 U1005 ( .A(n1131), .B(n1132), .Z(data_scrambled[9]) );
  IV U1006 ( .A(n1133), .Z(n1132) );
  OR2 U1007 ( .A(n1134), .B(data_66b_tpg[9]), .Z(n1133) );
  AN2 U1008 ( .A(data_66b_tpg[9]), .B(n1134), .Z(n1131) );
  AN2 U1009 ( .A(n1135), .B(n1136), .Z(n1134) );
  OR2 U1010 ( .A(n1137), .B(n[152]), .Z(n1136) );
  IV U1011 ( .A(n[133]), .Z(n1137) );
  OR2 U1012 ( .A(n1138), .B(n[133]), .Z(n1135) );
  OR2 U1013 ( .A(n1139), .B(n1140), .Z(data_scrambled[35]) );
  AN2 U1014 ( .A(n1141), .B(n1142), .Z(n1140) );
  IV U1015 ( .A(n1143), .Z(n1139) );
  OR2 U1016 ( .A(n1142), .B(n1141), .Z(n1143) );
  OR2 U1017 ( .A(n1144), .B(n1145), .Z(n1141) );
  AN2 U1018 ( .A(n[159]), .B(n890), .Z(n1145) );
  IV U1019 ( .A(n[178]), .Z(n890) );
  AN2 U1020 ( .A(n[178]), .B(n1146), .Z(n1144) );
  IV U1021 ( .A(data_66b_tpg[35]), .Z(n1142) );
  OR2 U1022 ( .A(n1147), .B(n1148), .Z(data_scrambled[34]) );
  AN2 U1023 ( .A(n1149), .B(n1150), .Z(n1148) );
  IV U1024 ( .A(n1151), .Z(n1147) );
  OR2 U1025 ( .A(n1150), .B(n1149), .Z(n1151) );
  OR2 U1026 ( .A(n1152), .B(n1153), .Z(n1149) );
  AN2 U1027 ( .A(n[158]), .B(n906), .Z(n1153) );
  IV U1028 ( .A(n[177]), .Z(n906) );
  AN2 U1029 ( .A(n[177]), .B(n898), .Z(n1152) );
  IV U1030 ( .A(n[158]), .Z(n898) );
  IV U1031 ( .A(data_66b_tpg[34]), .Z(n1150) );
  OR2 U1032 ( .A(n1154), .B(n1155), .Z(data_scrambled[33]) );
  AN2 U1033 ( .A(n1156), .B(n1157), .Z(n1155) );
  IV U1034 ( .A(n1158), .Z(n1154) );
  OR2 U1035 ( .A(n1157), .B(n1156), .Z(n1158) );
  OR2 U1036 ( .A(n1159), .B(n1160), .Z(n1156) );
  AN2 U1037 ( .A(n[157]), .B(n922), .Z(n1160) );
  IV U1038 ( .A(n[176]), .Z(n922) );
  AN2 U1039 ( .A(n[176]), .B(n914), .Z(n1159) );
  IV U1040 ( .A(n[157]), .Z(n914) );
  IV U1041 ( .A(data_66b_tpg[33]), .Z(n1157) );
  OR2 U1042 ( .A(n1161), .B(n1162), .Z(data_scrambled[32]) );
  AN2 U1043 ( .A(n1163), .B(n1164), .Z(n1162) );
  IV U1044 ( .A(n1165), .Z(n1161) );
  OR2 U1045 ( .A(n1164), .B(n1163), .Z(n1165) );
  OR2 U1046 ( .A(n1166), .B(n1167), .Z(n1163) );
  AN2 U1047 ( .A(n[156]), .B(n938), .Z(n1167) );
  IV U1048 ( .A(n[175]), .Z(n938) );
  AN2 U1049 ( .A(n[175]), .B(n930), .Z(n1166) );
  IV U1050 ( .A(n[156]), .Z(n930) );
  IV U1051 ( .A(data_66b_tpg[32]), .Z(n1164) );
  OR2 U1052 ( .A(n1168), .B(n1169), .Z(data_scrambled[31]) );
  AN2 U1053 ( .A(n1170), .B(n1171), .Z(n1169) );
  IV U1054 ( .A(n1172), .Z(n1168) );
  OR2 U1055 ( .A(n1171), .B(n1170), .Z(n1172) );
  OR2 U1056 ( .A(n1173), .B(n1174), .Z(n1170) );
  AN2 U1057 ( .A(n[155]), .B(n954), .Z(n1174) );
  IV U1058 ( .A(n[174]), .Z(n954) );
  AN2 U1059 ( .A(n[174]), .B(n946), .Z(n1173) );
  IV U1060 ( .A(n[155]), .Z(n946) );
  IV U1061 ( .A(data_66b_tpg[31]), .Z(n1171) );
  OR2 U1062 ( .A(n1175), .B(n1176), .Z(data_scrambled[30]) );
  AN2 U1063 ( .A(n1177), .B(n1178), .Z(n1176) );
  IV U1064 ( .A(n1179), .Z(n1175) );
  OR2 U1065 ( .A(n1178), .B(n1177), .Z(n1179) );
  OR2 U1066 ( .A(n1180), .B(n1181), .Z(n1177) );
  AN2 U1067 ( .A(n[154]), .B(n970), .Z(n1181) );
  IV U1068 ( .A(n[173]), .Z(n970) );
  AN2 U1069 ( .A(n[173]), .B(n962), .Z(n1180) );
  IV U1070 ( .A(n[154]), .Z(n962) );
  IV U1071 ( .A(data_66b_tpg[30]), .Z(n1178) );
  OR2 U1072 ( .A(n1182), .B(n1183), .Z(data_scrambled[29]) );
  AN2 U1073 ( .A(n1184), .B(n1185), .Z(n1183) );
  IV U1074 ( .A(n1186), .Z(n1182) );
  OR2 U1075 ( .A(n1185), .B(n1184), .Z(n1186) );
  OR2 U1076 ( .A(n1187), .B(n1188), .Z(n1184) );
  AN2 U1077 ( .A(n[153]), .B(n978), .Z(n1188) );
  IV U1078 ( .A(n[172]), .Z(n978) );
  AN2 U1079 ( .A(n[172]), .B(n1002), .Z(n1187) );
  IV U1080 ( .A(n[153]), .Z(n1002) );
  IV U1081 ( .A(data_66b_tpg[29]), .Z(n1185) );
  OR2 U1082 ( .A(n1189), .B(n1190), .Z(data_scrambled[28]) );
  AN2 U1083 ( .A(n1191), .B(n1192), .Z(n1190) );
  IV U1084 ( .A(n1193), .Z(n1189) );
  OR2 U1085 ( .A(n1192), .B(n1191), .Z(n1193) );
  OR2 U1086 ( .A(n1194), .B(n1195), .Z(n1191) );
  AN2 U1087 ( .A(n[152]), .B(n986), .Z(n1195) );
  IV U1088 ( .A(n[171]), .Z(n986) );
  AN2 U1089 ( .A(n[171]), .B(n1138), .Z(n1194) );
  IV U1090 ( .A(n[152]), .Z(n1138) );
  IV U1091 ( .A(data_66b_tpg[28]), .Z(n1192) );
  OR2 U1092 ( .A(n1196), .B(n1197), .Z(data_scrambled[27]) );
  AN2 U1093 ( .A(n1198), .B(n1199), .Z(n1197) );
  IV U1094 ( .A(n1200), .Z(n1196) );
  OR2 U1095 ( .A(n1199), .B(n1198), .Z(n1200) );
  OR2 U1096 ( .A(n1201), .B(n1202), .Z(n1198) );
  AN2 U1097 ( .A(n[151]), .B(n994), .Z(n1202) );
  IV U1098 ( .A(n[170]), .Z(n994) );
  AN2 U1099 ( .A(n[170]), .B(n1203), .Z(n1201) );
  IV U1100 ( .A(data_66b_tpg[27]), .Z(n1199) );
  OR2 U1101 ( .A(n1204), .B(n1205), .Z(data_scrambled[26]) );
  AN2 U1102 ( .A(n1206), .B(n1207), .Z(n1205) );
  IV U1103 ( .A(n1208), .Z(n1204) );
  OR2 U1104 ( .A(n1207), .B(n1206), .Z(n1208) );
  OR2 U1105 ( .A(n1209), .B(n1210), .Z(n1206) );
  AN2 U1106 ( .A(n[150]), .B(n1010), .Z(n1210) );
  IV U1107 ( .A(n[169]), .Z(n1010) );
  AN2 U1108 ( .A(n[169]), .B(n1211), .Z(n1209) );
  IV U1109 ( .A(data_66b_tpg[26]), .Z(n1207) );
  OR2 U1110 ( .A(n1212), .B(n1213), .Z(data_scrambled[8]) );
  IV U1111 ( .A(n1214), .Z(n1213) );
  OR2 U1112 ( .A(n1215), .B(data_66b_tpg[8]), .Z(n1214) );
  AN2 U1113 ( .A(data_66b_tpg[8]), .B(n1215), .Z(n1212) );
  AN2 U1114 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR2 U1115 ( .A(n1218), .B(n[151]), .Z(n1217) );
  IV U1116 ( .A(n[132]), .Z(n1218) );
  OR2 U1117 ( .A(n1203), .B(n[132]), .Z(n1216) );
  IV U1118 ( .A(n[151]), .Z(n1203) );
  OR2 U1119 ( .A(n1219), .B(n1220), .Z(data_scrambled[25]) );
  AN2 U1120 ( .A(n1221), .B(n1222), .Z(n1220) );
  IV U1121 ( .A(n1223), .Z(n1219) );
  OR2 U1122 ( .A(n1222), .B(n1221), .Z(n1223) );
  OR2 U1123 ( .A(n1224), .B(n1225), .Z(n1221) );
  AN2 U1124 ( .A(n[149]), .B(n1018), .Z(n1225) );
  IV U1125 ( .A(n[168]), .Z(n1018) );
  AN2 U1126 ( .A(n[168]), .B(n1226), .Z(n1224) );
  IV U1127 ( .A(data_66b_tpg[25]), .Z(n1222) );
  AN2 U1128 ( .A(n1227), .B(n1228), .Z(data_scrambled[24]) );
  OR2 U1129 ( .A(n1229), .B(n[148]), .Z(n1228) );
  IV U1130 ( .A(n1230), .Z(n1229) );
  OR2 U1131 ( .A(n1026), .B(n1230), .Z(n1227) );
  OR2 U1132 ( .A(n1231), .B(n1232), .Z(n1230) );
  AN2 U1133 ( .A(n[167]), .B(n1233), .Z(n1232) );
  IV U1134 ( .A(n483), .Z(n1233) );
  AN2 U1135 ( .A(n483), .B(n1034), .Z(n1231) );
  IV U1136 ( .A(n[167]), .Z(n1034) );
  IV U1137 ( .A(n[148]), .Z(n1026) );
  AN2 U1138 ( .A(n1234), .B(n1235), .Z(data_scrambled[23]) );
  OR2 U1139 ( .A(n1236), .B(n[147]), .Z(n1235) );
  IV U1140 ( .A(n1237), .Z(n1236) );
  OR2 U1141 ( .A(n1042), .B(n1237), .Z(n1234) );
  OR2 U1142 ( .A(n1238), .B(n1239), .Z(n1237) );
  AN2 U1143 ( .A(n[166]), .B(n1240), .Z(n1239) );
  IV U1144 ( .A(n484), .Z(n1240) );
  AN2 U1145 ( .A(n484), .B(n1050), .Z(n1238) );
  IV U1146 ( .A(n[166]), .Z(n1050) );
  IV U1147 ( .A(n[147]), .Z(n1042) );
  AN2 U1148 ( .A(n1241), .B(n1242), .Z(data_scrambled[22]) );
  OR2 U1149 ( .A(n1243), .B(n[146]), .Z(n1242) );
  IV U1150 ( .A(n1244), .Z(n1243) );
  OR2 U1151 ( .A(n1058), .B(n1244), .Z(n1241) );
  OR2 U1152 ( .A(n1245), .B(n1246), .Z(n1244) );
  AN2 U1153 ( .A(n[165]), .B(n1247), .Z(n1246) );
  IV U1154 ( .A(n485), .Z(n1247) );
  AN2 U1155 ( .A(n485), .B(n1066), .Z(n1245) );
  IV U1156 ( .A(n[165]), .Z(n1066) );
  IV U1157 ( .A(n[146]), .Z(n1058) );
  AN2 U1158 ( .A(n1248), .B(n1249), .Z(data_scrambled[21]) );
  OR2 U1159 ( .A(n1250), .B(n[145]), .Z(n1249) );
  IV U1160 ( .A(n1251), .Z(n1250) );
  OR2 U1161 ( .A(n1074), .B(n1251), .Z(n1248) );
  OR2 U1162 ( .A(n1252), .B(n1253), .Z(n1251) );
  AN2 U1163 ( .A(n[164]), .B(n1254), .Z(n1253) );
  IV U1164 ( .A(n486), .Z(n1254) );
  AN2 U1165 ( .A(n486), .B(n1082), .Z(n1252) );
  IV U1166 ( .A(n[164]), .Z(n1082) );
  IV U1167 ( .A(n[145]), .Z(n1074) );
  AN2 U1168 ( .A(n1255), .B(n1256), .Z(data_scrambled[20]) );
  OR2 U1169 ( .A(n1257), .B(n[144]), .Z(n1256) );
  IV U1170 ( .A(n1258), .Z(n1257) );
  OR2 U1171 ( .A(n1090), .B(n1258), .Z(n1255) );
  OR2 U1172 ( .A(n1259), .B(n1260), .Z(n1258) );
  AN2 U1173 ( .A(n[163]), .B(n1261), .Z(n1260) );
  IV U1174 ( .A(n487), .Z(n1261) );
  AN2 U1175 ( .A(n487), .B(n1098), .Z(n1259) );
  IV U1176 ( .A(n[163]), .Z(n1098) );
  IV U1177 ( .A(n[144]), .Z(n1090) );
  AN2 U1178 ( .A(n1262), .B(n1263), .Z(data_scrambled[19]) );
  OR2 U1179 ( .A(n1264), .B(n[143]), .Z(n1263) );
  IV U1180 ( .A(n1265), .Z(n1264) );
  OR2 U1181 ( .A(n1106), .B(n1265), .Z(n1262) );
  OR2 U1182 ( .A(n1266), .B(n1267), .Z(n1265) );
  AN2 U1183 ( .A(n[162]), .B(n1268), .Z(n1267) );
  IV U1184 ( .A(n488), .Z(n1268) );
  AN2 U1185 ( .A(n488), .B(n1114), .Z(n1266) );
  IV U1186 ( .A(n[162]), .Z(n1114) );
  IV U1187 ( .A(n[143]), .Z(n1106) );
  OR2 U1188 ( .A(n1269), .B(n1270), .Z(data_scrambled[18]) );
  IV U1189 ( .A(n1271), .Z(n1270) );
  OR2 U1190 ( .A(n1272), .B(data_66b_tpg[18]), .Z(n1271) );
  AN2 U1191 ( .A(data_66b_tpg[18]), .B(n1272), .Z(n1269) );
  AN2 U1192 ( .A(n1273), .B(n1274), .Z(n1272) );
  OR2 U1193 ( .A(n1275), .B(n[161]), .Z(n1274) );
  IV U1194 ( .A(n[142]), .Z(n1275) );
  OR2 U1195 ( .A(n1122), .B(n[142]), .Z(n1273) );
  IV U1196 ( .A(n[161]), .Z(n1122) );
  OR2 U1197 ( .A(n1276), .B(n1277), .Z(data_scrambled[17]) );
  IV U1198 ( .A(n1278), .Z(n1277) );
  OR2 U1199 ( .A(n1279), .B(data_66b_tpg[17]), .Z(n1278) );
  AN2 U1200 ( .A(data_66b_tpg[17]), .B(n1279), .Z(n1276) );
  AN2 U1201 ( .A(n1280), .B(n1281), .Z(n1279) );
  OR2 U1202 ( .A(n1282), .B(n[160]), .Z(n1281) );
  IV U1203 ( .A(n[141]), .Z(n1282) );
  OR2 U1204 ( .A(n1130), .B(n[141]), .Z(n1280) );
  IV U1205 ( .A(n[160]), .Z(n1130) );
  OR2 U1206 ( .A(n1283), .B(n1284), .Z(data_scrambled[16]) );
  IV U1207 ( .A(n1285), .Z(n1284) );
  OR2 U1208 ( .A(n1286), .B(data_66b_tpg[16]), .Z(n1285) );
  AN2 U1209 ( .A(data_66b_tpg[16]), .B(n1286), .Z(n1283) );
  AN2 U1210 ( .A(n1287), .B(n1288), .Z(n1286) );
  OR2 U1211 ( .A(n1289), .B(n[159]), .Z(n1288) );
  IV U1212 ( .A(n[140]), .Z(n1289) );
  OR2 U1213 ( .A(n1146), .B(n[140]), .Z(n1287) );
  IV U1214 ( .A(n[159]), .Z(n1146) );
  OR2 U1215 ( .A(n1290), .B(n1291), .Z(data_scrambled[7]) );
  IV U1216 ( .A(n1292), .Z(n1291) );
  OR2 U1217 ( .A(n1293), .B(data_66b_tpg[7]), .Z(n1292) );
  AN2 U1218 ( .A(data_66b_tpg[7]), .B(n1293), .Z(n1290) );
  AN2 U1219 ( .A(n1294), .B(n1295), .Z(n1293) );
  OR2 U1220 ( .A(n1296), .B(n[150]), .Z(n1295) );
  IV U1221 ( .A(n[131]), .Z(n1296) );
  OR2 U1222 ( .A(n1211), .B(n[131]), .Z(n1294) );
  IV U1223 ( .A(n[150]), .Z(n1211) );
  OR2 U1224 ( .A(n1297), .B(n1298), .Z(data_scrambled[6]) );
  IV U1225 ( .A(n1299), .Z(n1298) );
  OR2 U1226 ( .A(n1300), .B(data_66b_tpg[6]), .Z(n1299) );
  AN2 U1227 ( .A(data_66b_tpg[6]), .B(n1300), .Z(n1297) );
  AN2 U1228 ( .A(n1301), .B(n1302), .Z(n1300) );
  OR2 U1229 ( .A(n1303), .B(n[149]), .Z(n1302) );
  IV U1230 ( .A(n[130]), .Z(n1303) );
  OR2 U1231 ( .A(n1226), .B(n[130]), .Z(n1301) );
  IV U1232 ( .A(n[149]), .Z(n1226) );
endmodule

