// Benchmark "Huffman_jpeg_8" written by ABC on Fri Nov 21 18:10:47 2014

module Huffman_jpeg_8 ( clock, 
    in_0 , in_1 , in_2 , in_3 , in_4 , in_5 , in_6 , in_7 ,
    carestate, out  );
  input  clock;
  input  in_0 , in_1 , in_2 , in_3 , in_4 , in_5 , in_6 ,
    in_7 ;
  output carestate, out;
  reg reg_0 , reg_1 , reg_2 , reg_3 , reg_4 , reg_5 , reg_6 ,
    reg_7 , counter_0 , counter_1 , counter_2 , counter_3 ;
  wire n47_1, n56, n57_1, n58, n59, n60, n61, n62_1, n63, n64, n65, n66,
    n67_1, n72_1, n73, n74, n75, n76, n77_1, n78, n79, n80, n81, n83, n84,
    n22, n27, n32, n37, n42, n47, n52, n57, n62, n67, n72, n77;
  assign n47_1 = ~counter_0  & ~counter_1  & ~counter_2  & ~counter_3 ;
  assign n22 = n47_1 ? in_0  : reg_0 ;
  assign n27 = n47_1 ? in_1  : reg_1 ;
  assign n32 = n47_1 ? in_2  : reg_2 ;
  assign n37 = n47_1 ? in_3  : reg_3 ;
  assign n42 = n47_1 ? in_4  : reg_4 ;
  assign n47 = n47_1 ? in_5  : reg_5 ;
  assign n52 = n47_1 ? in_6  : reg_6 ;
  assign n57 = n47_1 ? in_7  : reg_7 ;
  assign n56 = ((in_4  ? (~in_5  & ~in_7 ) : (in_5  & in_7 )) & (in_0  | (~in_0  & in_6 ))) | (~in_5  & ((in_0  & ~in_4  & in_6 ) | (~in_0  & in_4  & ~in_6 ) | (in_0  & ~in_6  & in_7 ))) | (in_0  & ~in_4  & in_5  & ~in_7 ) | (~in_0  & in_1  & ~in_4  & ((~in_5  & in_6 ) | (in_5  & ~in_6 ) | (in_5  & in_6  & ~in_7 ))) | (~in_0  & ~in_1  & in_2  & ~in_4  & (in_6  ? (~in_5  ^ ~in_7 ) : in_5 )) | (in_3  & ~in_4  & ((~in_7  & ((in_2  & ~in_5  & (in_0  ? (in_1  & ~in_6 ) : (~in_1  & in_6 ))) | (~in_0  & ~in_1  & ~in_2  & in_5 ))) | (~in_0  & ~in_1  & ~in_2  & in_5  & ~in_6  & in_7 )));
  assign n57_1 = (~in_5  & (in_0  ? (in_4  ^ in_6 ) : (in_4  & ~in_6 ))) | (in_0  & ~in_4  & in_5 ) | (~in_0  & in_1  & ~in_4  & in_5 ) | (~in_5  & ((in_6  & ((in_4  & ~in_7 ) | (~in_0  & in_1  & ~in_4  & in_7 ))) | (~in_0  & in_1  & ~in_4  & ~in_6  & in_7 ))) | (~in_0  & ~in_1  & in_2  & ~in_4  & (in_5  ? (in_6  | (~in_6  & in_7 )) : (~in_6  & in_7 ))) | (~in_4  & ((~in_0  & ~in_1  & ((~in_7  & (in_2  ? (in_3  ? (in_5  & ~in_6 ) : (~in_5  & in_6 )) : (in_6  & (in_3  ^ in_5 )))) | (~in_2  & in_7  & (in_3  ? in_6  : (in_5  & ~in_6 ))))) | (in_0  & in_1  & in_2  & ~in_6  & in_7  & in_3  & ~in_5 )));
  assign n58 = ((in_4  ^ in_5 ) & ((in_0  & ~in_6  & in_7 ) | (~in_7  & (in_0  | (~in_0  & in_6 ))) | (~in_0  & in_1  & ~in_6 ))) | (~in_5  & ((in_0  & in_1  & ~in_4  & in_6 ) | (~in_0  & ~in_1  & in_4  & ~in_6 ) | (in_0  & ~in_1  & ~in_4  & in_6  & in_7 ))) | (~in_4  & in_5  & in_6  & in_7  & (in_0  | (~in_0  & in_1 ))) | (~in_0  & ~in_4  & ((in_6  & ((in_2  & (in_1  ? ~in_5  : (in_5  & in_7 ))) | (~in_5  & in_7  & ~in_1  & ~in_2 ))) | (~in_5  & ~in_6  & in_7  & in_1  & in_2 ))) | (~in_4  & ((~in_5  & ((in_2  & ((~in_1  & in_6  & (in_0  ? (in_3  & ~in_7 ) : (~in_3  ^ in_7 ))) | (in_0  & in_1  & ~in_6  & (~in_3  ^ ~in_7 )))) | (~in_0  & ~in_2  & ~in_6  & (in_1  ? (in_3  & in_7 ) : (~in_3  ^ in_7 ))))) | (~in_0  & ~in_1  & in_5  & ((~in_6  & (in_2  ? (~in_3  ^ in_7 ) : (~in_3  & ~in_7 ))) | (in_6  & in_7  & ~in_2  & in_3 )))));
  assign n59 = (~in_6  & (in_0  ? (in_4  ^ in_5 ) : (in_4  & ~in_5 ))) | (in_0  & ~in_4  & in_5  & in_6 ) | (in_1  & ~in_4  & (in_0  ? (~in_5  & in_6 ) : in_5 )) | (~in_5  & in_6  & (in_4  ? ~in_7  : (in_0  ? (~in_1  & in_7 ) : (in_1  & ~in_7 )))) | (~in_4  & ((in_7  & ((~in_2  & ~in_5  & (in_0  ? (in_1  & ~in_6 ) : (~in_1  ^ in_6 ))) | (~in_0  & ~in_1  & in_2  & in_5 ))) | (~in_0  & ~in_1  & in_2  & in_5  & ~in_7 ))) | (~in_4  & (in_0  ? (~in_5  & ((~in_1  & ((in_2  & (in_3  ? (~in_6  & in_7 ) : (in_6  & ~in_7 ))) | (in_6  & ~in_7  & ~in_2  & in_3 ))) | (in_1  & in_2  & in_3  & ~in_6  & ~in_7 ))) : ((~in_1  & ~in_2  & (in_3  ? (in_5  & in_7 ) : (~in_5  & ~in_7 ))) | (in_1  & in_2  & in_3  & ~in_5  & in_7 ) | (~in_3  & ((~in_1  & ((in_2  & ~in_5  & in_6 ) | (~in_2  & in_5  & ~in_6  & ~in_7 ))) | (~in_5  & ~in_6  & in_7  & in_1  & ~in_2 ))) | (~in_5  & ~in_6  & in_7  & ~in_1  & in_2  & in_3 ))));
  assign n60 = 1'b0;
  assign n61 = counter_3  | n60;
  assign n62_1 = counter_2  | n61;
  assign n63 = counter_1  | n62_1;
  assign n64 = counter_0  ^ ~n63;
  assign n65 = counter_1  ^ ~n62_1;
  assign n66 = counter_2  ^ ~n61;
  assign n67_1 = counter_3  ^ ~n60;
  assign n62 = n47_1 ? n56 : n64;
  assign n67 = n47_1 ? n57_1 : n65;
  assign n72 = n47_1 ? n58 : n66;
  assign n77 = n47_1 ? n59 : n67_1;
  assign n72_1 = in_0  ^ ~reg_0 ;
  assign n73 = in_1  ^ ~reg_1 ;
  assign n74 = in_2  ^ ~reg_2 ;
  assign n75 = in_3  ^ ~reg_3 ;
  assign n76 = in_4  ^ ~reg_4 ;
  assign n77_1 = in_5  ^ ~reg_5 ;
  assign n78 = in_6  ^ ~reg_6 ;
  assign n79 = in_7  ^ ~reg_7 ;
  assign n80 = n79 & n78 & n77_1 & n76 & n75 & n74 & n72_1 & n73;
  assign n81 = ((in_0  ^ in_1 ) & (in_5  ? in_4  : (in_4  ? (in_6  & in_7 ) : (~in_6  & ~in_7 )))) | (in_4  & (in_0  ^ ~in_1 ) & (in_5  | (~in_5  & in_6  & in_7 ))) | (~in_4  & ~in_5  & ~in_6  & ~in_7  & (in_0  ? (in_1  & ~in_2 ) : (~in_1  & in_2 ))) | (~in_4  & ~in_5  & ~in_6  & ~in_7  & ((~in_0  & ~in_1  & ~in_2  & in_3 ) | (in_0  & in_1  & in_2  & ~in_3 )));
  assign carestate = n47_1 ? ~n81 : n80;
  assign n83 = (in_6  & in_7 ) | (~in_6  & ~in_7 ) | ((in_6  ^ in_7 ) & ((~in_0  & ~in_1  & ~in_2  & in_3 ) | in_0  | (~in_0  & in_1 ) | (~in_0  & ~in_1  & in_2 ) | (~in_0  & ~in_1  & ~in_2  & ~in_3  & in_4 ) | (~in_0  & ~in_1  & ~in_2  & ~in_3  & ~in_4  & in_5 )));
  assign n84 = (~reg_4  & (((reg_5  ? (~reg_6  & ~reg_7 ) : (reg_6  & reg_7 )) & (reg_3  ? ((counter_1  & (counter_0  ? (reg_0  | (~counter_2  & ~reg_0  & reg_1 )) : ((reg_0  & reg_1  & counter_2  & ~counter_3 ) | (~counter_2  & counter_3  & ~reg_0  & ~reg_1 )))) | (counter_0  & ~counter_1  & (reg_0  | (~reg_0  & reg_1 )))) : (((counter_3  ? (~reg_0  & reg_1 ) : (reg_0  & ~reg_1 )) & ((counter_0  & counter_1  & ~counter_2 ) | (~counter_1  & (counter_0  | (~counter_0  & counter_2 ))))) | (reg_1  & ((~counter_0  & ~counter_1  & ~counter_2  & counter_3 ) | (counter_0  & ~counter_3  & (~counter_1  | (counter_1  & ~counter_2 ))) | (counter_0  & reg_0  & (counter_3  | (counter_1  & counter_2  & ~counter_3 ))))) | (counter_0  & reg_0  & ~reg_1  & (counter_3  | (counter_1  & counter_2  & ~counter_3 )))))) | (((reg_0  & (counter_2  ? ~reg_5  : (reg_1  & reg_5 ))) | (~counter_2  & ~reg_0  & reg_1  & ~reg_5 )) & ((~counter_0  & counter_1  & ~reg_6  & reg_7 ) | (counter_0  & ~counter_1  & reg_6  & ~reg_7 ))) | (reg_1  & ((counter_0  & ((reg_5  & (reg_7  | (counter_1  & reg_6  & ~reg_7 ) | (reg_6  & ~reg_7  & ~counter_1  & ~reg_0 ))) | (counter_1  & reg_0  & ~reg_5  & reg_6  & ~reg_7 ) | (~reg_7  & ((~counter_1  & reg_0  & reg_6  & (~counter_2  ^ reg_5 )) | (counter_1  & counter_2  & ~reg_0  & reg_5  & ~reg_6 ))) | (~counter_1  & ~counter_2  & reg_0  & ~reg_5  & ~reg_6  & reg_7 ))) | (~counter_0  & counter_1  & counter_2  & reg_6  & ~reg_7  & ~reg_0  & ~reg_5 ))) | (counter_0  & reg_0  & ~reg_1  & ((reg_5  & (reg_6  | (~reg_6  & reg_7 ))) | (~counter_1  & ~counter_2  & ~reg_5  & reg_6  & ~reg_7 ))) | (reg_7  & ((~counter_2  & ((~reg_1  & (counter_0  ? (~counter_1  & ~counter_3  & (reg_0  ? (~reg_5  & ~reg_6 ) : (reg_5  & reg_6 ))) : (counter_1  & counter_3  & reg_0  & (~reg_5  | (reg_5  & ~reg_6 ))))) | (~counter_0  & counter_1  & reg_1  & reg_5  & reg_6  & (~counter_3  ^ reg_0 )))) | (~counter_0  & counter_1  & counter_2  & reg_5  & (reg_0  | (~reg_0  & reg_1 )) & (~counter_3  ^ reg_6 )))) | (counter_1  & ~reg_7  & ((~counter_0  & ((reg_0  & ((reg_1  & ((~counter_2  & (counter_3  ? (reg_5  & ~reg_6 ) : (~reg_5  & reg_6 ))) | (counter_2  & counter_3  & reg_5  & reg_6 ))) | (counter_2  & ~reg_1  & (counter_3  ? reg_6  : (reg_5  & ~reg_6 ))))) | (~counter_2  & counter_3  & ~reg_0  & reg_6  & (~reg_1  ^ ~reg_5 )))) | (counter_0  & ~counter_2  & ~counter_3  & reg_0  & ~reg_1  & ~reg_5  & reg_6 ))) | (~counter_1  & ((reg_5  & ((~counter_2  & ~reg_1  & ((counter_0  & ~reg_0  & reg_3  & (~counter_3  ^ reg_7 )) | (~counter_0  & counter_3  & reg_0  & ~reg_3  & ~reg_7 ))) | (~counter_0  & counter_2  & ~counter_3  & ~reg_0  & reg_1  & ~reg_3  & ~reg_7 ) | (~reg_0  & ((reg_3  & ((reg_7  & (counter_0  ? (~reg_1  & (counter_2  ? reg_6  : (~counter_3  & ~reg_6 ))) : (counter_2  ? ((counter_3  ^ reg_1 ) & ~reg_6 ) : (counter_3  & reg_6 )))) | (~reg_1  & ~reg_7  & ((counter_0  & reg_6  & (counter_2  ^ counter_3 )) | (~counter_0  & counter_2  & counter_3  & ~reg_6 ))))) | (~counter_0  & counter_3  & ~reg_3  & ((reg_1  & (counter_2  ? (reg_6  ^ reg_7 ) : (~reg_6  & reg_7 ))) | (reg_6  & ~reg_7  & ~counter_2  & ~reg_1 ))))) | (~counter_0  & counter_3  & reg_0  & ((reg_1  & (counter_2  ? (reg_3  ? (~reg_6  & reg_7 ) : (reg_6  & ~reg_7 )) : (reg_3  ? (reg_6  & reg_7 ) : (reg_6  ^ reg_7 )))) | (~counter_2  & ~reg_1  & reg_7  & (~reg_3  ^ reg_6 )))))) | (~counter_0  & ~reg_5  & (counter_2  ? ((reg_3  & (reg_0  ? ((counter_3  & ~reg_1  & ~reg_6  & reg_7 ) | (~counter_3  & reg_1  & reg_6  & ~reg_7 )) : ((reg_6  & (counter_3  ? (~reg_1  ^ reg_7 ) : (~reg_1  & reg_7 ))) | (~reg_6  & reg_7  & ~counter_3  & ~reg_1 )))) | (~counter_3  & ~reg_0  & reg_1  & ~reg_3  & (reg_6  ^ reg_7 ))) : (counter_3  & ((reg_1  & ((~reg_0  & (reg_3  ? (reg_6  & ~reg_7 ) : (~reg_6  & reg_7 ))) | (reg_0  & ~reg_3  & reg_6  & ~reg_7 ))) | (reg_0  & ~reg_1  & reg_3  & reg_7 ))))))) | (counter_1  & (reg_0  ? ((~counter_0  & ((~counter_3  & ((~reg_3  & ((counter_2  & ~reg_7  & (reg_1  ? (reg_5  & ~reg_6 ) : (~reg_5  & reg_6 ))) | (~counter_2  & reg_1  & ~reg_5  & reg_6  & reg_7 ))) | (~counter_2  & reg_3  & ~reg_6  & reg_7  & (~reg_1  ^ ~reg_5 )))) | (~counter_2  & counter_3  & reg_1  & ~reg_6  & reg_7  & ~reg_3  & ~reg_5 ))) | (counter_3  & ~reg_1  & counter_0  & ~counter_2  & reg_6  & ~reg_7  & reg_3  & ~reg_5 )) : ((reg_5  & (counter_0  ? (~reg_1  & reg_3  & reg_6  & reg_7 ) : ((~reg_7  & (counter_2  ? ((~counter_3  & reg_1  & ~reg_3  & reg_6 ) | (counter_3  & ~reg_1  & reg_3  & ~reg_6 )) : ((~counter_3  & ~reg_1  & ~reg_3  & reg_6 ) | (reg_3  & ~reg_6  & counter_3  & reg_1 )))) | (~counter_2  & ~reg_1  & ~reg_3  & reg_7  & (~counter_3  ^ reg_6 ))))) | (~counter_0  & ~reg_5  & reg_7  & ((counter_2  & ((~counter_3  & reg_3  & (reg_1  ^ reg_6 )) | (~reg_3  & reg_6  & counter_3  & reg_1 ))) | (~counter_2  & ~counter_3  & reg_1  & reg_3  & reg_6 )))))))) | (reg_4  & ~reg_5  & ((~reg_7  & (((~reg_1  ^ reg_6 ) & (((~counter_2  ^ reg_3 ) & (counter_0  | (~counter_0  & counter_3  & reg_0 ))) | ((counter_2  ^ reg_3 ) & (counter_0  | (~counter_0  & counter_1  & counter_3  & reg_0 ))) | (~counter_0  & counter_1  & ~counter_2  & ~counter_3  & reg_0 ))) | (counter_3  & (reg_0  ? (((reg_1  ^ reg_6 ) & (counter_0  | (~counter_0  & counter_1  & counter_2 ) | (~counter_0  & ~counter_1  & ~counter_2  & ~reg_3 ))) | (~counter_0  & counter_1  & ~counter_2  & ~reg_1  & reg_6 )) : ((counter_1  & (counter_0  ? (reg_1  ^ reg_6 ) : reg_1 )) | (counter_0  & ~counter_1  & (reg_1  ^ reg_6 )) | (~counter_0  & ~counter_1  & (counter_2  ? (reg_1  ? (reg_3  & reg_6 ) : (~reg_3  & ~reg_6 )) : (reg_1  & ~reg_3 )))))) | (~counter_3  & ((counter_0  & ~counter_1  & (reg_1  ^ reg_6 )) | (counter_1  & (counter_0  ? (reg_1  ^ reg_6 ) : (((~reg_1  ^ reg_3 ) & (counter_2  ? reg_6  : (~reg_0  & ~reg_6 ))) | (counter_2  & (((~reg_1  ^ ~reg_3 ) & reg_6 ) | (reg_0  & reg_1  & reg_3  & ~reg_6 ))) | (~counter_2  & reg_0  & ~reg_1  & reg_3  & reg_6 )))))))) | (~reg_6  & reg_7  & ((counter_1  & counter_2  & ~counter_3  & reg_3 ) | (~counter_1  & ~counter_2  & counter_3  & ~reg_3 ) | (counter_0  & ((counter_1  & ~counter_2 ) | (~counter_1  & counter_2 ) | (counter_1  & counter_2  & counter_3 ) | (~counter_1  & ~counter_2  & ~counter_3 ) | (~counter_1  & ~counter_2  & counter_3  & reg_3 ) | (counter_1  & counter_2  & ~counter_3  & ~reg_3 ))) | (~counter_0  & counter_2  & reg_1  & (counter_1  ? (counter_3  | (~counter_3  & ~reg_3 )) : (counter_3  & ~reg_3 ))) | (~counter_0  & ((counter_1  & reg_0  & ((~reg_1  & ((counter_2  & counter_3 ) | (~counter_2  & ~counter_3 ) | (counter_2  & ~counter_3  & ~reg_3 ))) | (reg_1  & ~reg_3  & ~counter_2  & ~counter_3 ))) | (~counter_1  & counter_2  & ~counter_3  & ~reg_0  & ~reg_1  & ~reg_3 ))))))) | (reg_2  & ((~reg_0  & (counter_1  ? ((~reg_1  & ((~counter_2  & ((reg_3  & ((~reg_4  & reg_5  & (counter_0  ? ~reg_7  : (~counter_3  & reg_7 ))) | (~counter_0  & counter_3  & reg_4  & ~reg_5  & ~reg_7 ))) | (counter_0  & ~reg_3  & ~reg_4  & reg_5  & reg_7 ))) | (~counter_0  & counter_2  & counter_3  & ~reg_5  & ~reg_7  & reg_3  & reg_4 ))) | (~counter_0  & ~counter_2  & counter_3  & reg_1  & reg_5  & ~reg_7  & ~reg_3  & ~reg_4 )) : (counter_2  ? (counter_0  ? (~reg_1  & ~reg_4  & reg_5  & (~reg_3  | (counter_3  & reg_3  & ~reg_7 ))) : ((~reg_4  & ((counter_3  & reg_5  & (reg_1  ? (reg_3  & reg_7 ) : (~reg_3  & ~reg_7 ))) | (~counter_3  & ~reg_1  & ~reg_3  & ~reg_5  & reg_7 ))) | (~counter_3  & reg_3  & reg_4  & ~reg_5  & ~reg_7 ))) : (~reg_1  & ~reg_3  & ~reg_4  & ((counter_3  & (counter_0  ? reg_5  : (~reg_5  & reg_7 ))) | (counter_0  & ~counter_3  & reg_5  & ~reg_7 )))))) | (~counter_0  & counter_2  & reg_0  & ((~counter_1  & ((reg_1  & ((~reg_3  & ~reg_4  & ((reg_7  & (counter_3  | (~counter_3  & ~reg_5 ))) | (~counter_3  & reg_5  & ~reg_7 ))) | (~counter_3  & reg_3  & reg_4  & ~reg_5  & ~reg_7 ))) | (reg_4  & ~reg_5  & ~reg_7  & ~counter_3  & ~reg_1  & reg_3 ))) | (counter_1  & ~counter_3  & reg_1  & ~reg_5  & ~reg_7  & reg_3  & ~reg_4 ))))) | (~counter_0  & ~reg_2  & ((~reg_4  & ((reg_5  & ((~reg_1  & (counter_1  ? (~reg_0  & reg_3  & (counter_2  ? (~counter_3  & ~reg_7 ) : (counter_3  & reg_7 ))) : (counter_2  & reg_0  & ~reg_3  & reg_7 ))) | (~counter_1  & counter_2  & ~counter_3  & reg_0  & reg_1  & (~reg_3  ^ ~reg_7 )))) | (~counter_1  & counter_2  & reg_0  & ~reg_5  & reg_7  & (counter_3  ? (~reg_1  & ~reg_3 ) : (reg_1  & reg_3 ))))) | (~counter_1  & reg_4  & ~reg_5  & ~reg_7  & ((counter_2  & ~counter_3  & ~reg_3  & (reg_0  | (~reg_0  & reg_1 ))) | (~counter_2  & counter_3  & ~reg_0  & ~reg_1  & reg_3 ))))) | (~counter_0  & ((~reg_5  & (counter_3  ? ((reg_2  & ((reg_3  & ((~counter_1  & ~reg_6  & ((counter_2  & ~reg_0  & ~reg_1  & reg_4 ) | (~counter_2  & reg_0  & reg_1  & ~reg_4 ))) | (counter_1  & counter_2  & ~reg_0  & ~reg_1  & ~reg_4  & reg_6 ))) | (counter_1  & ~reg_0  & ~reg_1  & ~reg_3  & ~reg_4  & reg_6 ))) | (counter_1  & ~counter_2  & ~reg_0  & ~reg_1  & ~reg_2  & ~reg_3  & reg_4  & ~reg_6 ) | (~counter_2  & (((reg_2  ? (reg_3  & reg_7 ) : (~reg_3  & ~reg_7 )) & ((~counter_1  & ~reg_0  & ~reg_1  & ~reg_4  & reg_6 ) | (counter_1  & reg_0  & reg_1  & reg_4  & ~reg_6 ))) | (reg_6  & (reg_0  ? (~reg_4  & ((counter_1  & reg_1  & (reg_2  ? (reg_3  ^ ~reg_7 ) : (~reg_3  ^ ~reg_7 ))) | (reg_2  & ~reg_3  & ~reg_7  & ~counter_1  & ~reg_1 ))) : ((reg_1  & ~reg_2  & reg_3  & ~reg_4  & reg_7 ) | (~reg_1  & reg_2  & ~reg_3  & reg_4  & ~reg_7 ) | (counter_1  & ~reg_4  & ((reg_1  & ~reg_2  & ~reg_3  & reg_7 ) | (~reg_1  & reg_2  & reg_3  & ~reg_7 )))))) | (reg_3  & ~reg_4  & ~reg_6  & ((counter_1  & ((reg_0  & reg_1  & (reg_2  ^ reg_7 )) | (~reg_0  & ~reg_1  & reg_2  & reg_7 ))) | (~counter_1  & ~reg_0  & reg_1  & reg_2  & reg_7 ))))) | (counter_2  & (reg_2  ? (reg_3  ? ((~reg_6  & ((reg_7  & (reg_1  ^ reg_4 ) & (counter_1  ^ reg_0 )) | (counter_1  & reg_0  & reg_1  & ~reg_4  & ~reg_7 ))) | (~counter_1  & ~reg_4  & reg_6  & ((~reg_7  & (reg_0  | (~reg_0  & reg_1 ))) | (~reg_0  & ~reg_1  & reg_7 )))) : ((reg_4  & ((~reg_0  & ((counter_1  & ~reg_1  & (reg_6  ^ reg_7 )) | (reg_6  & ~reg_7  & ~counter_1  & reg_1 ))) | (~counter_1  & reg_0  & ~reg_7  & (~reg_1  ^ reg_6 )))) | (~counter_1  & ~reg_0  & ~reg_1  & ~reg_4  & reg_6  & reg_7 ))) : ((~reg_0  & ((~counter_1  & ((reg_4  & ((~reg_6  & (reg_1  ? (reg_3  ^ ~reg_7 ) : (~reg_3  & reg_7 ))) | (~reg_1  & reg_3  & reg_6  & ~reg_7 ))) | (~reg_3  & ~reg_4  & ~reg_7  & (~reg_1  ^ reg_6 )))) | (~reg_4  & reg_6  & reg_7  & counter_1  & reg_1  & reg_3 ))) | (~counter_1  & reg_0  & ((~reg_3  & ~reg_7  & (reg_1  ? (reg_4  ^ reg_6 ) : reg_6 )) | (reg_1  & reg_3  & reg_4  & ~reg_6  & reg_7 ))))))) : (reg_4  ? (((reg_0  ? (reg_2  & ~reg_3 ) : (~reg_2  & reg_3 )) & ((~counter_1  & counter_2  & ~reg_6  & reg_7 ) | (counter_1  & ~counter_2  & ~reg_1  & reg_6  & ~reg_7 ))) | (~reg_6  & ((counter_2  & ((reg_7  & ((~counter_1  & ((reg_0  & ~reg_2  & reg_3 ) | (reg_2  & ~reg_3  & ~reg_0  & reg_1 ))) | (counter_1  & ~reg_0  & ~reg_1  & reg_2  & ~reg_3 ))) | (counter_1  & ~reg_7  & ((~reg_0  & ~reg_1  & (reg_2  ^ reg_3 )) | (reg_2  & ~reg_3  & reg_0  & reg_1 ))))) | (counter_1  & ~counter_2  & ((reg_1  & (reg_0  ^ reg_2 ) & (reg_3  ^ ~reg_7 )) | (~reg_0  & ~reg_1  & ~reg_2  & ~reg_3  & reg_7 )))))) : (reg_6  ? ((counter_2  & ((reg_3  & ((~reg_1  & ((~reg_7  & (counter_1  ? (reg_0  ^ reg_2 ) : (~reg_0  & reg_2 ))) | (~counter_1  & reg_0  & reg_2  & reg_7 ))) | (~counter_1  & ~reg_0  & reg_1  & ~reg_2  & reg_7 ))) | (reg_2  & ~reg_3  & ((reg_0  & reg_1  & (~counter_1  ^ reg_7 )) | (counter_1  & ~reg_0  & ~reg_1 ))))) | (counter_1  & ~counter_2  & ((~reg_2  & (reg_1  ? (reg_0  ? (reg_3  & reg_7 ) : (~reg_3  ^ ~reg_7 )) : (~reg_0  ^ ~reg_3 ))) | (~reg_0  & ~reg_1  & reg_2  & ~reg_3  & ~reg_7 )))) : ((reg_0  & ((reg_7  & ((counter_1  & ~counter_2  & ~reg_3  & (reg_1  ^ reg_2 )) | (~reg_1  & ~reg_2  & reg_3  & ~counter_1  & counter_2 ))) | (~counter_1  & counter_2  & reg_1  & reg_2  & reg_3  & ~reg_7 ))) | (counter_1  & ~reg_0  & reg_2  & reg_7  & (counter_2  ? (reg_1  & ~reg_3 ) : ~reg_1 ))))))) | (~reg_4  & reg_5  & (((reg_2  ^ reg_3 ) & ((~reg_0  & ((counter_1  & ((counter_2  & counter_3  & ~reg_1  & ~reg_6  & reg_7 ) | (~counter_2  & ~counter_3  & reg_1  & reg_6  & ~reg_7 ))) | (reg_1  & reg_6  & ~reg_7  & ~counter_1  & ~counter_2  & counter_3 ))) | (~counter_1  & counter_2  & reg_0  & ~reg_1  & ~reg_7  & (~counter_3  ^ ~reg_6 )))) | ((reg_2  ^ reg_6 ) & ((~counter_3  & ((counter_2  & ((~counter_1  & reg_0  & reg_3  & reg_7 ) | (~reg_1  & ~reg_3  & ~reg_7  & counter_1  & ~reg_0 ))) | (counter_1  & ~counter_2  & ~reg_1  & (reg_0  ? (~reg_3  & reg_7 ) : (reg_3  & ~reg_7 ))))) | (~counter_1  & counter_2  & counter_3  & reg_0  & reg_1  & reg_3  & ~reg_7 ))) | (reg_3  & (reg_6  ? (counter_1  ? (counter_2  ? (~reg_0  & ((counter_3  & ~reg_1  & reg_2  & reg_7 ) | (~reg_7  & (counter_3  ? (~reg_1  ^ reg_2 ) : (reg_1  & ~reg_2 ))))) : (reg_0  & ((~counter_3  & (reg_1  ? (reg_2  & ~reg_7 ) : (~reg_2  & reg_7 ))) | (counter_3  & ~reg_1  & reg_2  & reg_7 )))) : (counter_2  & ((reg_7  & ((counter_3  & (reg_0  ? (~reg_1  ^ reg_2 ) : (~reg_1  & ~reg_2 ))) | (reg_1  & ~reg_2  & ~counter_3  & ~reg_0 ))) | (counter_3  & ~reg_1  & reg_2  & ~reg_7 )))) : ((~reg_0  & (reg_1  ? ((~reg_2  & ((~counter_1  & (counter_2  ? ~reg_7  : (counter_3  & reg_7 ))) | (counter_1  & ~counter_2  & ~counter_3  & reg_7 ))) | (counter_1  & ~counter_2  & reg_2  & (~counter_3  ^ reg_7 ))) : ((~counter_1  & ((counter_2  & ~counter_3  & reg_2 ) | (~counter_2  & counter_3  & ~reg_2  & ~reg_7 ))) | (counter_1  & counter_2  & ~counter_3  & ~reg_2  & reg_7 )))) | (counter_1  & ~counter_2  & ~counter_3  & reg_0  & ~reg_1  & reg_2  & ~reg_7 )))) | (~reg_3  & ((~reg_0  & (reg_6  ? (reg_7  & ((~reg_2  & (counter_1  ? (~reg_1  & (counter_2  | (~counter_2  & ~counter_3 ))) : (counter_2  ? (~counter_3  & reg_1 ) : (counter_3  & ~reg_1 )))) | (~counter_1  & counter_2  & counter_3  & reg_1  & reg_2 ))) : (((counter_3  ? (reg_2  & reg_7 ) : (~reg_2  & ~reg_7 )) & (counter_1  ? (~counter_2  & reg_1 ) : (counter_2  & ~reg_1 ))) | (~reg_1  & (counter_1  ? (counter_3  & reg_2  & (~counter_2  | (counter_2  & ~reg_7 ))) : (~reg_2  & (counter_2  ? (~counter_3  & reg_7 ) : (counter_3  & ~reg_7 )))))))) | (counter_1  & ~counter_2  & counter_3  & reg_0  & ~reg_1  & reg_2  & reg_6  & reg_7 ))))))) | (counter_0  & reg_2  & ~reg_4  & ((~reg_5  & (reg_0  ? (reg_3  ? ((~counter_3  & (counter_1  ? ((~counter_2  & reg_1  & ~reg_6  & reg_7 ) | (reg_6  & ~reg_7  & counter_2  & ~reg_1 )) : (reg_1  & ~reg_6  & (counter_2  | (~counter_2  & ~reg_7 ))))) | (~counter_1  & counter_3  & ~reg_6  & ((reg_1  & (counter_2  | (~counter_2  & ~reg_7 ))) | (~counter_2  & ~reg_1  & reg_7 )))) : ((~counter_1  & counter_2  & ~counter_3  & reg_1  & ~reg_6  & reg_7 ) | (~reg_1  & reg_6  & ~reg_7  & counter_1  & ~counter_2  & counter_3 ))) : (reg_6  & ((~counter_1  & (counter_2  ? (reg_1  & ~reg_7 ) : (~reg_1  & reg_7 ))) | (counter_1  & counter_2  & ~counter_3  & reg_1  & reg_7 ) | (reg_3  & ((~counter_1  & ~counter_3  & ~reg_1  & (counter_2  ^ ~reg_7 )) | (counter_1  & counter_2  & counter_3  & reg_1  & reg_7 ))))))) | (~reg_0  & ~reg_1  & reg_5  & (((counter_3  ? (reg_3  & ~reg_7 ) : (~reg_3  & reg_7 )) & (counter_1  ? (counter_2  & reg_6 ) : (~counter_2  & ~reg_6 ))) | (counter_2  & ((~reg_3  & reg_6  & counter_1  & counter_3 ) | (reg_3  & ~reg_6  & ~counter_1  & ~counter_3 ) | (reg_3  & ((~reg_6  & reg_7  & (counter_1  | (~counter_1  & counter_3 ))) | (reg_6  & ~reg_7  & counter_1  & ~counter_3 ))) | (~reg_3  & reg_6  & ~reg_7  & counter_1  & ~counter_3 ))) | (counter_1  & ~counter_2  & (reg_3  ? (~reg_6  & reg_7 ) : (reg_6  & ~reg_7 )))))));
  assign out = n47_1 ? n83 : n84;
  always @ (posedge clock) begin
    reg_0  <= n22;
    reg_1  <= n27;
    reg_2  <= n32;
    reg_3  <= n37;
    reg_4  <= n42;
    reg_5  <= n47;
    reg_6  <= n52;
    reg_7  <= n57;
    counter_0  <= n62;
    counter_1  <= n67;
    counter_2  <= n72;
    counter_3  <= n77;
  end
  initial begin
    reg_0  <= 1'b0;
    reg_1  <= 1'b0;
    reg_2  <= 1'b0;
    reg_3  <= 1'b0;
    reg_4  <= 1'b0;
    reg_5  <= 1'b0;
    reg_6  <= 1'b0;
    reg_7  <= 1'b0;
    counter_0  <= 1'b0;
    counter_1  <= 1'b0;
    counter_2  <= 1'b0;
    counter_3  <= 1'b0;
  end
endmodule


