
module XGXSSYNTH_ENC_8B10B ( bad_code, bad_disp, clk, encode_data_in, konstant, 
        rst, disp_out, encode_data_out, assertion_shengyushen );
  input [7:0] encode_data_in;
  output [9:0] encode_data_out;
  input bad_code, bad_disp, clk, konstant, rst;
  output disp_out, assertion_shengyushen;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n12, n13, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n140, n141, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n182, n183, n188, n189, n190,
         n191, n194, n195, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n216, n221,
         n224, n226, n233, n240, n241, n242, n243, n244, n258, n259, U5_Z_0,
         U5_DATA1_0, U4_Z_0, n297, n302, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n352, n353, n354,
         n355, n356, n357, n358, n359, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431;
  wire   [187:184] n;

  OR2 C692 ( .A(n203), .B(bad_code), .Z(encode_data_out[0]) );
  AN2 C690 ( .A(n202), .B(n1), .Z(encode_data_out[1]) );
  OR2 C689 ( .A(n201), .B(bad_code), .Z(encode_data_out[2]) );
  OR2 C688 ( .A(n200), .B(bad_code), .Z(encode_data_out[3]) );
  OR2 C687 ( .A(n199), .B(bad_code), .Z(encode_data_out[4]) );
  OR2 C686 ( .A(n198), .B(bad_code), .Z(encode_data_out[5]) );
  AN2 C684 ( .A(n207), .B(n1), .Z(encode_data_out[6]) );
  OR2 C683 ( .A(n206), .B(bad_code), .Z(encode_data_out[7]) );
  AN2 C681 ( .A(n205), .B(n1), .Z(encode_data_out[8]) );
  IV I_50 ( .A(bad_code), .Z(n1) );
  AN2 C679 ( .A(n204), .B(n1), .Z(encode_data_out[9]) );
  OR2 C674 ( .A(n306), .B(n179), .Z(n3) );
  AN2 C673 ( .A(n191), .B(n3), .Z(n2) );
  OR2 C672 ( .A(n180), .B(n182), .Z(n5) );
  AN2 C670 ( .A(n312), .B(n5), .Z(n4) );
  OR2 C669 ( .A(n4), .B(n2), .Z(n178) );
  AN2 C666 ( .A(n183), .B(n190), .Z(n7) );
  AN2 C665 ( .A(n7), .B(n6), .Z(n182) );
  AN2 C662 ( .A(n6), .B(n310), .Z(n8) );
  OR2 C661 ( .A(n8), .B(n188), .Z(n[184]) );
  OR2 C660 ( .A(n194), .B(n308), .Z(n[186]) );
  AN2 C658 ( .A(n195), .B(n302), .Z(n[187]) );
  AN2 C657 ( .A(n189), .B(n100), .Z(n188) );
  AN2 C655 ( .A(n312), .B(n90), .Z(n13) );
  AN2 C654 ( .A(n191), .B(n311), .Z(n15) );
  OR2 C653 ( .A(n15), .B(n13), .Z(n12) );
  OR2 C652 ( .A(n12), .B(n190), .Z(n189) );
  IV I_46 ( .A(rst), .Z(n216) );
  OR2 C635 ( .A(n221), .B(n136), .Z(n16) );
  OR2 C632 ( .A(n97), .B(n95), .Z(n221) );
  OR2 C629 ( .A(n233), .B(n226), .Z(n17) );
  IV I_44 ( .A(n258), .Z(n19) );
  AN2 C626 ( .A(n19), .B(konstant), .Z(n18) );
  OR2 C625 ( .A(n102), .B(n226), .Z(n22) );
  AN2 C624 ( .A(U5_Z_0), .B(n22), .Z(n21) );
  AN2 C622 ( .A(n297), .B(n233), .Z(n23) );
  OR2 C621 ( .A(n23), .B(n21), .Z(n20) );
  OR2 C620 ( .A(n20), .B(n18), .Z(n214) );
  AN2 C619 ( .A(n93), .B(konstant), .Z(n25) );
  OR2 C618 ( .A(n73), .B(n71), .Z(n30) );
  OR2 C617 ( .A(n30), .B(n67), .Z(n29) );
  OR2 C616 ( .A(n29), .B(n63), .Z(n28) );
  OR2 C615 ( .A(n28), .B(n59), .Z(n27) );
  OR2 C614 ( .A(n27), .B(n58), .Z(n26) );
  OR2 C613 ( .A(n26), .B(n25), .Z(n226) );
  OR2 C606 ( .A(n88), .B(n86), .Z(n35) );
  OR2 C605 ( .A(n35), .B(n84), .Z(n34) );
  OR2 C604 ( .A(n34), .B(n82), .Z(n33) );
  OR2 C603 ( .A(n33), .B(n80), .Z(n32) );
  OR2 C602 ( .A(n32), .B(n77), .Z(n31) );
  OR2 C601 ( .A(n31), .B(n75), .Z(n233) );
  AN2 C594 ( .A(n93), .B(konstant), .Z(n36) );
  AN2 C590 ( .A(n44), .B(n43), .Z(n42) );
  AN2 C589 ( .A(n42), .B(n176), .Z(n41) );
  AN2 C587 ( .A(n113), .B(n46), .Z(n45) );
  OR2 C586 ( .A(n45), .B(n41), .Z(n40) );
  OR2 C585 ( .A(n40), .B(n109), .Z(n39) );
  OR2 C584 ( .A(n39), .B(n107), .Z(n38) );
  OR2 C583 ( .A(n38), .B(n58), .Z(n37) );
  OR2 C582 ( .A(n37), .B(n36), .Z(n240) );
  OR2 C581 ( .A(n123), .B(n118), .Z(n48) );
  OR2 C580 ( .A(n48), .B(n115), .Z(n47) );
  OR2 C578 ( .A(n49), .B(n47), .Z(n241) );
  AN2 C576 ( .A(encode_data_in[3]), .B(n52), .Z(n242) );
  OR2 C575 ( .A(encode_data_in[2]), .B(n132), .Z(n50) );
  OR2 C574 ( .A(n50), .B(n75), .Z(n243) );
  IV I_42 ( .A(n130), .Z(n52) );
  AN2 C572 ( .A(encode_data_in[1]), .B(n52), .Z(n51) );
  OR2 C571 ( .A(n51), .B(n132), .Z(n244) );
  OR2 C558 ( .A(n93), .B(n259), .Z(n258) );
  OR2 C557 ( .A(n71), .B(n67), .Z(n54) );
  OR2 C556 ( .A(n54), .B(n63), .Z(n53) );
  OR2 C555 ( .A(n53), .B(n59), .Z(n259) );
  OR2 C553 ( .A(n166), .B(n156), .Z(n57) );
  OR2 C552 ( .A(n57), .B(n147), .Z(n56) );
  AN2 C551 ( .A(konstant), .B(n56), .Z(n55) );
  OR2 C550 ( .A(n177), .B(n55), .Z(assertion_shengyushen) );
  AN2 C501 ( .A(encode_data_in[4]), .B(n130), .Z(n58) );
  IV I_41 ( .A(n60), .Z(n59) );
  OR2 C496 ( .A(n176), .B(n61), .Z(n60) );
  OR2 C495 ( .A(n175), .B(n62), .Z(n61) );
  OR2 C494 ( .A(n174), .B(n121), .Z(n62) );
  IV I_40 ( .A(n64), .Z(n63) );
  OR2 C487 ( .A(n176), .B(n65), .Z(n64) );
  OR2 C486 ( .A(n175), .B(n66), .Z(n65) );
  OR2 C485 ( .A(n174), .B(n126), .Z(n66) );
  IV I_39 ( .A(n68), .Z(n67) );
  OR2 C478 ( .A(n176), .B(n69), .Z(n68) );
  OR2 C477 ( .A(n175), .B(n70), .Z(n69) );
  OR2 C476 ( .A(encode_data_in[2]), .B(n106), .Z(n70) );
  IV I_38 ( .A(n72), .Z(n71) );
  OR2 C469 ( .A(n176), .B(n104), .Z(n72) );
  IV I_37 ( .A(n74), .Z(n73) );
  OR2 C460 ( .A(n176), .B(n133), .Z(n74) );
  IV I_36 ( .A(n76), .Z(n75) );
  OR2 C454 ( .A(n176), .B(n129), .Z(n76) );
  IV I_35 ( .A(n78), .Z(n77) );
  OR2 C447 ( .A(encode_data_in[4]), .B(n79), .Z(n78) );
  OR2 C446 ( .A(n175), .B(n105), .Z(n79) );
  IV I_34 ( .A(n81), .Z(n80) );
  OR2 C438 ( .A(encode_data_in[4]), .B(n129), .Z(n81) );
  IV I_33 ( .A(n83), .Z(n82) );
  OR2 C432 ( .A(encode_data_in[4]), .B(n116), .Z(n83) );
  IV I_32 ( .A(n85), .Z(n84) );
  OR2 C426 ( .A(encode_data_in[4]), .B(n119), .Z(n85) );
  IV I_31 ( .A(n87), .Z(n86) );
  OR2 C420 ( .A(encode_data_in[4]), .B(n124), .Z(n87) );
  IV I_30 ( .A(n89), .Z(n88) );
  OR2 C414 ( .A(encode_data_in[4]), .B(n133), .Z(n89) );
  AN2 C410 ( .A(n198), .B(n199), .Z(n90) );
  OR2 C408 ( .A(n198), .B(n199), .Z(n92) );
  IV I_28 ( .A(n94), .Z(n93) );
  OR2 C406 ( .A(n176), .B(n111), .Z(n94) );
  IV I_27 ( .A(n96), .Z(n95) );
  OR2 C398 ( .A(n155), .B(n99), .Z(n96) );
  IV I_26 ( .A(n98), .Z(n97) );
  OR2 C394 ( .A(encode_data_in[7]), .B(n99), .Z(n98) );
  OR2 C393 ( .A(encode_data_in[6]), .B(encode_data_in[5]), .Z(n99) );
  AN2 C392 ( .A(n[185]), .B(n101), .Z(n100) );
  AN2 C391 ( .A(n194), .B(n195), .Z(n101) );
  IV I_25 ( .A(n103), .Z(n102) );
  OR2 C389 ( .A(encode_data_in[4]), .B(n104), .Z(n103) );
  OR2 C388 ( .A(encode_data_in[3]), .B(n105), .Z(n104) );
  OR2 C387 ( .A(n174), .B(n106), .Z(n105) );
  OR2 C386 ( .A(n122), .B(n127), .Z(n106) );
  IV I_24 ( .A(n108), .Z(n107) );
  OR2 C381 ( .A(n176), .B(n116), .Z(n108) );
  IV I_23 ( .A(n110), .Z(n109) );
  OR2 C374 ( .A(encode_data_in[4]), .B(n111), .Z(n110) );
  OR2 C373 ( .A(n175), .B(n117), .Z(n111) );
  AN2 C368 ( .A(encode_data_in[1]), .B(encode_data_in[0]), .Z(n112) );
  IV I_22 ( .A(n114), .Z(n113) );
  OR2 C366 ( .A(encode_data_in[3]), .B(encode_data_in[2]), .Z(n114) );
  IV I_21 ( .A(n116), .Z(n115) );
  OR2 C364 ( .A(encode_data_in[3]), .B(n117), .Z(n116) );
  OR2 C363 ( .A(n174), .B(n135), .Z(n117) );
  IV I_20 ( .A(n119), .Z(n118) );
  OR2 C359 ( .A(encode_data_in[3]), .B(n120), .Z(n119) );
  OR2 C358 ( .A(encode_data_in[2]), .B(n121), .Z(n120) );
  OR2 C357 ( .A(n122), .B(encode_data_in[0]), .Z(n121) );
  IV I_19 ( .A(encode_data_in[1]), .Z(n122) );
  IV I_18 ( .A(n124), .Z(n123) );
  OR2 C354 ( .A(encode_data_in[3]), .B(n125), .Z(n124) );
  OR2 C353 ( .A(encode_data_in[2]), .B(n126), .Z(n125) );
  OR2 C352 ( .A(encode_data_in[1]), .B(n127), .Z(n126) );
  IV I_17 ( .A(encode_data_in[0]), .Z(n127) );
  IV I_16 ( .A(n129), .Z(n128) );
  OR2 C349 ( .A(n175), .B(n134), .Z(n129) );
  AN2 C345 ( .A(encode_data_in[3]), .B(n131), .Z(n130) );
  AN2 C344 ( .A(encode_data_in[2]), .B(n112), .Z(n131) );
  IV I_15 ( .A(n133), .Z(n132) );
  OR2 C341 ( .A(encode_data_in[3]), .B(n134), .Z(n133) );
  OR2 C340 ( .A(encode_data_in[2]), .B(n135), .Z(n134) );
  OR2 C339 ( .A(encode_data_in[1]), .B(encode_data_in[0]), .Z(n135) );
  AN2 C338 ( .A(encode_data_in[7]), .B(n137), .Z(n136) );
  AN2 C337 ( .A(encode_data_in[6]), .B(encode_data_in[5]), .Z(n137) );
  IV I_14 ( .A(bad_disp), .Z(n138) );
  OR2 C334 ( .A(n[185]), .B(n141), .Z(n140) );
  OR2 C333 ( .A(n309), .B(n307), .Z(n141) );
  OR2 C329 ( .A(n[185]), .B(n146), .Z(n145) );
  OR2 C328 ( .A(n194), .B(n195), .Z(n146) );
  IV I_9 ( .A(n148), .Z(n147) );
  OR2 C326 ( .A(encode_data_in[0]), .B(n149), .Z(n148) );
  OR2 C325 ( .A(encode_data_in[1]), .B(n150), .Z(n149) );
  OR2 C324 ( .A(n174), .B(n151), .Z(n150) );
  OR2 C323 ( .A(n175), .B(n152), .Z(n151) );
  OR2 C322 ( .A(n176), .B(n153), .Z(n152) );
  OR2 C321 ( .A(n164), .B(n154), .Z(n153) );
  OR2 C320 ( .A(encode_data_in[6]), .B(n155), .Z(n154) );
  IV I_8 ( .A(encode_data_in[7]), .Z(n155) );
  IV I_7 ( .A(n157), .Z(n156) );
  OR2 C313 ( .A(encode_data_in[0]), .B(n158), .Z(n157) );
  OR2 C312 ( .A(encode_data_in[1]), .B(n159), .Z(n158) );
  OR2 C311 ( .A(n174), .B(n160), .Z(n159) );
  OR2 C310 ( .A(n175), .B(n161), .Z(n160) );
  OR2 C309 ( .A(n176), .B(n162), .Z(n161) );
  OR2 C308 ( .A(n164), .B(n163), .Z(n162) );
  OR2 C307 ( .A(n165), .B(encode_data_in[7]), .Z(n163) );
  IV I_6 ( .A(encode_data_in[5]), .Z(n164) );
  IV I_5 ( .A(encode_data_in[6]), .Z(n165) );
  IV I_4 ( .A(n167), .Z(n166) );
  OR2 C300 ( .A(encode_data_in[0]), .B(n168), .Z(n167) );
  OR2 C299 ( .A(encode_data_in[1]), .B(n169), .Z(n168) );
  OR2 C298 ( .A(n174), .B(n170), .Z(n169) );
  OR2 C297 ( .A(n175), .B(n171), .Z(n170) );
  OR2 C296 ( .A(n176), .B(n172), .Z(n171) );
  OR2 C295 ( .A(encode_data_in[5]), .B(n173), .Z(n172) );
  OR2 C294 ( .A(encode_data_in[6]), .B(encode_data_in[7]), .Z(n173) );
  IV I_3 ( .A(encode_data_in[2]), .Z(n174) );
  IV I_2 ( .A(encode_data_in[3]), .Z(n175) );
  IV I_1 ( .A(encode_data_in[4]), .Z(n176) );
  IV I_0 ( .A(konstant), .Z(n177) );
  FD1 disp_lat_reg ( .D(U4_Z_0), .CP(clk), .Q(U5_DATA1_0) );
  FD1 konstant_latch_reg ( .D(konstant), .CP(clk), .Q(n190) );
  FD1 ip_data_latch_reg_2_ ( .D(encode_data_in[5]), .CP(clk), .Q(n195) );
  FD1 ip_data_latch_reg_1_ ( .D(encode_data_in[6]), .CP(clk), .Q(n194) );
  FD1 ip_data_latch_reg_0_ ( .D(encode_data_in[7]), .CP(clk), .Q(n[185]) );
  FD1 disp_lat_fix_latch_reg ( .D(U5_Z_0), .CP(clk), .Q(disp_out) );
  FD1 data_out_latch_reg_5_ ( .D(n213), .CP(clk), .Q(n203) );
  FD1 data_out_latch_reg_4_ ( .D(n212), .CP(clk), .Q(n202) );
  FD1 data_out_latch_reg_3_ ( .D(n211), .CP(clk), .Q(n201) );
  FD1 data_out_latch_reg_2_ ( .D(n210), .CP(clk), .Q(n200) );
  FD1 data_out_latch_reg_1_ ( .D(n209), .CP(clk), .Q(n199) );
  FD1 data_out_latch_reg_0_ ( .D(n208), .CP(clk), .Q(n198) );
  FD1 kx_latch_reg ( .D(n93), .CP(clk), .Q(n183) );
  FD1 plus34_latch_reg ( .D(n221), .CP(clk), .Q(n180) );
  FD1 minus34b_latch_reg ( .D(n136), .CP(clk), .Q(n179) );
  FD1 i_disp_latch_reg ( .D(n224), .CP(clk), .Q(n191) );
  IV U25 ( .A(n355), .Z(n313) );
  IV U26 ( .A(n353), .Z(n314) );
  IV U27 ( .A(encode_data_in[4]), .Z(n315) );
  IV U28 ( .A(encode_data_in[3]), .Z(n316) );
  IV U29 ( .A(encode_data_in[2]), .Z(n317) );
  IV U30 ( .A(n357), .Z(n318) );
  IV U31 ( .A(encode_data_in[0]), .Z(n319) );
  OR2 U32 ( .A(n352), .B(n314), .Z(n49) );
  OR2 U33 ( .A(n315), .B(n128), .Z(n353) );
  AN2 U34 ( .A(n128), .B(n315), .Z(n352) );
  OR2 U35 ( .A(n354), .B(n313), .Z(n46) );
  OR2 U36 ( .A(n315), .B(n112), .Z(n355) );
  AN2 U37 ( .A(n112), .B(n315), .Z(n354) );
  OR2 U38 ( .A(n356), .B(n318), .Z(n44) );
  OR2 U39 ( .A(n319), .B(encode_data_in[1]), .Z(n357) );
  AN2 U40 ( .A(encode_data_in[1]), .B(n319), .Z(n356) );
  OR2 U41 ( .A(n358), .B(n359), .Z(n43) );
  AN2 U42 ( .A(encode_data_in[2]), .B(n316), .Z(n359) );
  AN2 U43 ( .A(encode_data_in[3]), .B(n317), .Z(n358) );
  OR2 U87 ( .A(n389), .B(n390), .Z(n6) );
  AN2 U88 ( .A(n194), .B(n307), .Z(n390) );
  AN2 U89 ( .A(n195), .B(n309), .Z(n389) );
  IV U90 ( .A(n191), .Z(n312) );
  IV U91 ( .A(n92), .Z(n311) );
  IV U92 ( .A(n194), .Z(n309) );
  IV U93 ( .A(n145), .Z(n308) );
  IV U94 ( .A(n195), .Z(n307) );
  IV U95 ( .A(n140), .Z(n306) );
  IV U96 ( .A(n188), .Z(n302) );
  OR2 U97 ( .A(n391), .B(n392), .Z(n213) );
  AN2 U98 ( .A(n319), .B(n214), .Z(n392) );
  AN2 U99 ( .A(encode_data_in[0]), .B(n393), .Z(n391) );
  OR2 U100 ( .A(n394), .B(n395), .Z(n212) );
  AN2 U101 ( .A(n214), .B(n396), .Z(n395) );
  IV U102 ( .A(n244), .Z(n396) );
  AN2 U103 ( .A(n244), .B(n393), .Z(n394) );
  OR2 U104 ( .A(n397), .B(n398), .Z(n211) );
  AN2 U105 ( .A(n214), .B(n399), .Z(n398) );
  IV U106 ( .A(n243), .Z(n399) );
  AN2 U107 ( .A(n243), .B(n393), .Z(n397) );
  OR2 U108 ( .A(n400), .B(n401), .Z(n210) );
  AN2 U109 ( .A(n214), .B(n402), .Z(n401) );
  IV U110 ( .A(n242), .Z(n402) );
  AN2 U111 ( .A(n242), .B(n393), .Z(n400) );
  OR2 U112 ( .A(n403), .B(n404), .Z(n209) );
  AN2 U113 ( .A(n214), .B(n405), .Z(n404) );
  IV U114 ( .A(n241), .Z(n405) );
  AN2 U115 ( .A(n241), .B(n393), .Z(n403) );
  OR2 U116 ( .A(n406), .B(n407), .Z(n208) );
  AN2 U117 ( .A(n214), .B(n408), .Z(n407) );
  IV U118 ( .A(n240), .Z(n408) );
  AN2 U119 ( .A(n240), .B(n393), .Z(n406) );
  IV U120 ( .A(n214), .Z(n393) );
  OR2 U121 ( .A(n409), .B(n410), .Z(n207) );
  AN2 U122 ( .A(n178), .B(n411), .Z(n410) );
  IV U123 ( .A(n[187]), .Z(n411) );
  AN2 U124 ( .A(n[187]), .B(n412), .Z(n409) );
  OR2 U125 ( .A(n413), .B(n414), .Z(n206) );
  AN2 U126 ( .A(n178), .B(n415), .Z(n414) );
  IV U127 ( .A(n[186]), .Z(n415) );
  AN2 U128 ( .A(n[186]), .B(n412), .Z(n413) );
  OR2 U129 ( .A(n416), .B(n417), .Z(n205) );
  AN2 U130 ( .A(n178), .B(n310), .Z(n417) );
  IV U131 ( .A(n[185]), .Z(n310) );
  AN2 U132 ( .A(n[185]), .B(n412), .Z(n416) );
  OR2 U133 ( .A(n418), .B(n419), .Z(n204) );
  AN2 U134 ( .A(n178), .B(n420), .Z(n419) );
  IV U135 ( .A(n[184]), .Z(n420) );
  AN2 U136 ( .A(n[184]), .B(n412), .Z(n418) );
  IV U137 ( .A(n178), .Z(n412) );
  AN2 U138 ( .A(n216), .B(n421), .Z(U4_Z_0) );
  OR2 U139 ( .A(n422), .B(n423), .Z(n421) );
  AN2 U140 ( .A(n224), .B(n424), .Z(n423) );
  IV U141 ( .A(n16), .Z(n424) );
  IV U142 ( .A(n425), .Z(n224) );
  AN2 U143 ( .A(n16), .B(n425), .Z(n422) );
  AN2 U144 ( .A(n426), .B(n427), .Z(n425) );
  OR2 U145 ( .A(n297), .B(n17), .Z(n427) );
  IV U146 ( .A(U5_Z_0), .Z(n297) );
  OR2 U147 ( .A(n428), .B(U5_Z_0), .Z(n426) );
  OR2 U148 ( .A(n429), .B(n430), .Z(U5_Z_0) );
  AN2 U149 ( .A(n138), .B(U5_DATA1_0), .Z(n430) );
  AN2 U150 ( .A(bad_disp), .B(n431), .Z(n429) );
  IV U151 ( .A(U5_DATA1_0), .Z(n431) );
  IV U152 ( .A(n17), .Z(n428) );
endmodule

