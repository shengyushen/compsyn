
module scrambler ( CLK, reset, data_66b_tpg, data_scrambled, 
        assertion_shengyushen );
  input [63:0] data_66b_tpg;
  output [63:0] data_scrambled;
  input CLK, reset;
  output assertion_shengyushen;
  wire   U4_DATA2_0, U4_DATA2_2, U4_DATA2_3, U4_DATA2_4, U4_DATA2_5,
         U4_DATA2_8, U4_DATA2_9, U4_DATA2_10, U4_DATA2_11, U4_DATA2_12, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n479, n480, n481, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n654, n656, n657, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691;
  wire   [167:124] n;

  FDS2P data_prev_reg_56_ ( .CR(data_scrambled[62]), .D(n504), .CP(CLK), .Q(
        n489), .QN(n654) );
  FDS2P data_prev_reg_36_ ( .CR(n661), .D(data_scrambled[42]), .CP(CLK), .Q(
        n[160]), .QN(n622) );
  FDS2P data_prev_reg_25_ ( .CR(n659), .D(data_scrambled[31]), .CP(CLK), .Q(
        n[149]), .QN(n579) );
  FDS2P data_prev_reg_29_ ( .CR(n656), .D(data_scrambled[35]), .CP(CLK), .Q(
        n[153]), .QN(n587) );
  FDS2P data_prev_reg_40_ ( .CR(n502), .D(data_scrambled[46]), .CP(CLK), .Q(
        n608), .QN(n488) );
  FDS2P data_prev_reg_34_ ( .CR(n662), .D(data_scrambled[40]), .CP(CLK), .Q(
        n607), .QN(n498) );
  FDS2P data_prev_reg_37_ ( .CR(n500), .D(data_scrambled[43]), .CP(CLK), .Q(
        n606), .QN(n496) );
  FDS2P data_prev_reg_39_ ( .CR(assertion_shengyushen), .D(data_scrambled[45]), 
        .CP(CLK), .Q(n605), .QN(n487) );
  FDS2P data_prev_reg_33_ ( .CR(n503), .D(data_scrambled[39]), .CP(CLK), .Q(
        n[157]), .QN(n591) );
  FDS2P data_prev_reg_30_ ( .CR(n501), .D(data_scrambled[36]), .CP(CLK), .Q(
        n604), .QN(n494) );
  FDS2P data_prev_reg_28_ ( .CR(n659), .D(data_scrambled[34]), .CP(CLK), .Q(
        n603), .QN(n492) );
  FDS2P data_prev_reg_35_ ( .CR(n656), .D(data_scrambled[41]), .CP(CLK), .Q(
        n602), .QN(n490) );
  FDS2 data_prev_reg_14_ ( .CR(n701), .D(data_scrambled[20]), .CP(CLK), .Q(
        n[138]), .QN() );
  FDS2 data_prev_reg_7_ ( .CR(assertion_shengyushen), .D(data_scrambled[13]), 
        .CP(CLK), .Q(n[131]), .QN() );
  FDS2 data_prev_reg_6_ ( .CR(n501), .D(data_scrambled[12]), .CP(CLK), .Q(
        n[130]), .QN() );
  FDS2 data_prev_reg_1_ ( .CR(assertion_shengyushen), .D(data_scrambled[7]), 
        .CP(CLK), .Q(n[125]), .QN() );
  FDS2 data_prev_reg_3_ ( .CR(n502), .D(data_scrambled[9]), .CP(CLK), .Q(
        n[127]), .QN() );
  FDS2 data_prev_reg_10_ ( .CR(n575), .D(U4_DATA2_10), .CP(CLK), .Q(n[134]), 
        .QN() );
  FDS2 data_prev_reg_18_ ( .CR(n503), .D(data_scrambled[24]), .CP(CLK), .Q(
        n[142]), .QN() );
  FDS2 data_prev_reg_17_ ( .CR(data_scrambled[23]), .D(n575), .CP(CLK), .Q(
        n[141]), .QN() );
  FDS2 data_prev_reg_16_ ( .CR(data_scrambled[22]), .D(n575), .CP(CLK), .Q(
        n[140]), .QN() );
  FDS2 data_prev_reg_15_ ( .CR(n501), .D(data_scrambled[21]), .CP(CLK), .Q(
        n[139]), .QN() );
  FDS2 data_prev_reg_13_ ( .CR(n503), .D(data_scrambled[19]), .CP(CLK), .Q(
        n[137]), .QN() );
  FDS2 data_prev_reg_12_ ( .CR(n502), .D(U4_DATA2_12), .CP(CLK), .Q(n[136]), 
        .QN() );
  FDS2 data_prev_reg_5_ ( .CR(n503), .D(U4_DATA2_5), .CP(CLK), .Q(n[129]), 
        .QN() );
  FDS2 data_prev_reg_0_ ( .CR(n656), .D(U4_DATA2_0), .CP(CLK), .Q(n[124]), 
        .QN() );
  FDS2 data_prev_reg_9_ ( .CR(n501), .D(data_scrambled[15]), .CP(CLK), .Q(
        n[133]), .QN() );
  FDS2 data_prev_reg_4_ ( .CR(n504), .D(data_scrambled[10]), .CP(CLK), .Q(
        n[128]), .QN() );
  FDS2 data_prev_reg_11_ ( .CR(n501), .D(data_scrambled[17]), .CP(CLK), .Q(
        n[135]), .QN() );
  FDS2 data_prev_reg_2_ ( .CR(n503), .D(data_scrambled[8]), .CP(CLK), .Q(
        n[126]), .QN() );
  FDS2 data_prev_reg_46_ ( .CR(data_scrambled[52]), .D(n504), .CP(CLK), .Q(
        n552), .QN(n472) );
  FDS2 data_prev_reg_48_ ( .CR(data_scrambled[54]), .D(n501), .CP(CLK), .Q(
        n553), .QN(n474) );
  FDS2 data_prev_reg_52_ ( .CR(data_scrambled[58]), .D(n503), .CP(CLK), .Q(
        n554), .QN(n476) );
  FDS2 data_prev_reg_51_ ( .CR(data_scrambled[57]), .D(n502), .CP(CLK), .Q(
        n555), .QN(n468) );
  FDS2P data_prev_reg_49_ ( .CR(n502), .D(data_scrambled[55]), .CP(CLK), .Q(
        n613), .QN() );
  FDS2P data_prev_reg_45_ ( .CR(data_scrambled[51]), .D(n659), .CP(CLK), .Q(
        n486), .QN(n508) );
  FDS2P data_prev_reg_53_ ( .CR(data_scrambled[59]), .D(n504), .CP(CLK), .Q(
        n611), .QN() );
  FDS2P data_prev_reg_47_ ( .CR(data_scrambled[53]), .D(n662), .CP(CLK), .Q(
        n610), .QN() );
  FDS2P data_prev_reg_57_ ( .CR(data_scrambled[63]), .D(n503), .CP(CLK), .Q(
        n485), .QN(n506) );
  FDS2P data_prev_reg_50_ ( .CR(data_scrambled[56]), .D(n659), .CP(CLK), .Q(
        n484), .QN(n505) );
  FDS2P data_prev_reg_54_ ( .CR(data_scrambled[60]), .D(n501), .CP(CLK), .Q(
        n612), .QN() );
  FDS2P data_prev_reg_44_ ( .CR(data_scrambled[50]), .D(n504), .CP(CLK), .Q(
        n609), .QN(n470) );
  FDS2P data_prev_reg_55_ ( .CR(data_scrambled[61]), .D(n502), .CP(CLK), .Q(
        n483), .QN(n507) );
  FDS2P data_prev_reg_27_ ( .CR(data_scrambled[33]), .D(assertion_shengyushen), 
        .CP(CLK), .Q(n[151]), .QN(n583) );
  FDS2P data_prev_reg_23_ ( .CR(data_scrambled[29]), .D(n656), .CP(CLK), .Q(
        n[147]), .QN() );
  FDS2P data_prev_reg_21_ ( .CR(data_scrambled[27]), .D(n502), .CP(CLK), .Q(
        n[145]), .QN() );
  FDS2P data_prev_reg_24_ ( .CR(data_scrambled[30]), .D(n503), .CP(CLK), .Q(
        n[148]), .QN() );
  FDS2P data_prev_reg_22_ ( .CR(data_scrambled[28]), .D(n504), .CP(CLK), .Q(
        n[146]), .QN() );
  FDS2P data_prev_reg_19_ ( .CR(data_scrambled[25]), .D(n701), .CP(CLK), .Q(
        n[143]), .QN() );
  FDS2P data_prev_reg_20_ ( .CR(data_scrambled[26]), .D(n504), .CP(CLK), .Q(
        n[144]), .QN() );
  FDS2P data_prev_reg_43_ ( .CR(data_scrambled[49]), .D(n502), .CP(CLK), .Q(
        n[167]), .QN() );
  FDS2P data_prev_reg_8_ ( .CR(U4_DATA2_8), .D(n502), .CP(CLK), .Q(n[132]), 
        .QN() );
  FDS2P data_prev_reg_38_ ( .CR(data_scrambled[44]), .D(n661), .CP(CLK), .Q(
        n[162]), .QN(n626) );
  FDS2P data_prev_reg_42_ ( .CR(data_scrambled[48]), .D(n501), .CP(CLK), .Q(
        n[166]), .QN(n618) );
  FDS2P data_prev_reg_41_ ( .CR(data_scrambled[47]), .D(n504), .CP(CLK), .Q(
        n[165]), .QN(n634) );
  FDS2P data_prev_reg_31_ ( .CR(data_scrambled[37]), .D(n501), .CP(CLK), .Q(), 
        .QN(n573) );
  FDS2P data_prev_reg_32_ ( .CR(data_scrambled[38]), .D(n503), .CP(CLK), .Q(), 
        .QN(n569) );
  FDS2P data_prev_reg_26_ ( .CR(data_scrambled[32]), .D(n701), .CP(CLK), .Q(), 
        .QN(n571) );
  EN U157 ( .A(n[125]), .B(data_66b_tpg[1]), .Z(n671) );
  B2I U158 ( .A(n610), .Z1(), .Z2(n556) );
  B2I U159 ( .A(n613), .Z1(), .Z2(n559) );
  EN U160 ( .A(n[133]), .B(data_66b_tpg[9]), .Z(n669) );
  IVP U161 ( .A(data_scrambled[2]), .Z(n687) );
  B2I U162 ( .A(n611), .Z1(), .Z2(n557) );
  B2I U163 ( .A(n612), .Z1(), .Z2(n558) );
  IVP U164 ( .A(n535), .Z(n689) );
  IVDA U165 ( .A(n627), .Y(), .Z(n566) );
  IVDA U166 ( .A(n623), .Y(), .Z(n565) );
  IVDA U167 ( .A(n630), .Y(), .Z(n567) );
  IVP U168 ( .A(n556), .Z(n537) );
  IVP U169 ( .A(n559), .Z(n540) );
  EO U170 ( .A(n679), .B(n574), .Z(n515) );
  EO U171 ( .A(n680), .B(n570), .Z(n513) );
  IVP U172 ( .A(n557), .Z(n538) );
  IVDA U173 ( .A(n619), .Y(), .Z(n564) );
  EO U174 ( .A(n664), .B(n572), .Z(n514) );
  IVP U175 ( .A(n558), .Z(n539) );
  IVDA U176 ( .A(n635), .Y(), .Z(n568) );
  EO U177 ( .A(n[147]), .B(n674), .Z(n699) );
  EN U178 ( .A(data_66b_tpg[59]), .B(n640), .Z(data_scrambled[59]) );
  IVDA U179 ( .A(n692), .Y(data_scrambled[24]), .Z(n479) );
  EN U180 ( .A(n[126]), .B(data_66b_tpg[2]), .Z(n672) );
  IVP U181 ( .A(n609), .Z(n471) );
  EO U182 ( .A(n603), .B(data_66b_tpg[28]), .Z(n432) );
  EN U183 ( .A(n432), .B(n537), .Z(data_scrambled[28]) );
  EO U184 ( .A(n537), .B(data_66b_tpg[47]), .Z(n433) );
  EN U185 ( .A(n433), .B(data_scrambled[8]), .Z(data_scrambled[47]) );
  ND2 U186 ( .A(n484), .B(n510), .Z(n434) );
  ND2 U187 ( .A(n434), .B(n524), .Z(n435) );
  EO U188 ( .A(n435), .B(data_66b_tpg[50]), .Z(data_scrambled[50]) );
  ND2 U189 ( .A(n542), .B(n616), .Z(n436) );
  ND2 U190 ( .A(n436), .B(n615), .Z(n437) );
  EO U191 ( .A(n437), .B(data_66b_tpg[48]), .Z(data_scrambled[48]) );
  EO U192 ( .A(n540), .B(data_66b_tpg[49]), .Z(n438) );
  EN U193 ( .A(n438), .B(data_scrambled[10]), .Z(data_scrambled[49]) );
  EN U194 ( .A(data_scrambled[17]), .B(data_66b_tpg[56]), .Z(n439) );
  EN U195 ( .A(n439), .B(n489), .Z(data_scrambled[56]) );
  EO U196 ( .A(n538), .B(data_66b_tpg[53]), .Z(n440) );
  EN U197 ( .A(n440), .B(data_scrambled[14]), .Z(data_scrambled[53]) );
  ND2 U198 ( .A(n544), .B(n515), .Z(n441) );
  ND2 U199 ( .A(n441), .B(n639), .Z(n442) );
  EO U200 ( .A(n442), .B(data_66b_tpg[51]), .Z(data_scrambled[51]) );
  ND2 U201 ( .A(data_scrambled[19]), .B(n480), .Z(n443) );
  ND2 U202 ( .A(n443), .B(n545), .Z(n444) );
  EO U203 ( .A(n444), .B(data_66b_tpg[58]), .Z(data_scrambled[58]) );
  EO U204 ( .A(n606), .B(data_66b_tpg[37]), .Z(n445) );
  EN U205 ( .A(n445), .B(n481), .Z(data_scrambled[37]) );
  EO U206 ( .A(n604), .B(data_66b_tpg[30]), .Z(n446) );
  EN U207 ( .A(n446), .B(n540), .Z(data_scrambled[30]) );
  ND2 U208 ( .A(n535), .B(n548), .Z(n447) );
  ND2 U209 ( .A(n447), .B(n547), .Z(n448) );
  EO U210 ( .A(n448), .B(data_66b_tpg[61]), .Z(data_scrambled[61]) );
  ND2 U211 ( .A(n485), .B(n511), .Z(n449) );
  ND2 U212 ( .A(n449), .B(n528), .Z(n450) );
  EO U213 ( .A(n450), .B(data_66b_tpg[57]), .Z(data_scrambled[57]) );
  EO U214 ( .A(n539), .B(data_66b_tpg[54]), .Z(n451) );
  EN U215 ( .A(n451), .B(data_scrambled[15]), .Z(data_scrambled[54]) );
  ND2 U216 ( .A(n543), .B(n513), .Z(n452) );
  ND2 U217 ( .A(n452), .B(n638), .Z(n453) );
  EO U218 ( .A(n453), .B(data_66b_tpg[52]), .Z(data_scrambled[52]) );
  ND2 U219 ( .A(data_scrambled[2]), .B(n634), .Z(n454) );
  ND2 U220 ( .A(n454), .B(n633), .Z(n455) );
  EO U221 ( .A(n455), .B(data_66b_tpg[41]), .Z(data_scrambled[41]) );
  EO U222 ( .A(n607), .B(data_66b_tpg[34]), .Z(n456) );
  EN U223 ( .A(n456), .B(n538), .Z(data_scrambled[34]) );
  ND2 U224 ( .A(n486), .B(n509), .Z(n457) );
  ND2 U225 ( .A(n457), .B(n523), .Z(n458) );
  EO U226 ( .A(n458), .B(data_66b_tpg[45]), .Z(data_scrambled[45]) );
  EO U227 ( .A(n566), .B(data_66b_tpg[32]), .Z(data_scrambled[32]) );
  EO U228 ( .A(n565), .B(data_66b_tpg[38]), .Z(data_scrambled[38]) );
  EO U229 ( .A(n567), .B(data_66b_tpg[26]), .Z(data_scrambled[26]) );
  EO U230 ( .A(n479), .B(data_66b_tpg[63]), .Z(n459) );
  EN U231 ( .A(n459), .B(data_scrambled[5]), .Z(data_scrambled[63]) );
  EO U232 ( .A(n564), .B(data_66b_tpg[36]), .Z(data_scrambled[36]) );
  ND2 U233 ( .A(n605), .B(n480), .Z(n460) );
  ND2 U234 ( .A(n460), .B(n592), .Z(n461) );
  EO U235 ( .A(n461), .B(data_66b_tpg[39]), .Z(data_scrambled[39]) );
  EO U236 ( .A(n532), .B(data_66b_tpg[43]), .Z(n462) );
  EN U237 ( .A(n462), .B(n660), .Z(data_scrambled[43]) );
  ND2 U238 ( .A(n541), .B(n514), .Z(n463) );
  ND2 U239 ( .A(n463), .B(n614), .Z(n464) );
  EO U240 ( .A(n464), .B(data_66b_tpg[46]), .Z(data_scrambled[46]) );
  EO U241 ( .A(n602), .B(data_66b_tpg[35]), .Z(n465) );
  EN U242 ( .A(n465), .B(n539), .Z(data_scrambled[35]) );
  EO U243 ( .A(n568), .B(data_66b_tpg[31]), .Z(data_scrambled[31]) );
  ND2 U244 ( .A(n535), .B(n618), .Z(n466) );
  ND2 U245 ( .A(n466), .B(n617), .Z(n467) );
  EO U246 ( .A(n467), .B(data_66b_tpg[42]), .Z(data_scrambled[42]) );
  B4I U247 ( .A(n529), .Z(n570) );
  IVP U248 ( .A(reset), .Z(n575) );
  EO U249 ( .A(n691), .B(data_66b_tpg[24]), .Z(n692) );
  B4I U250 ( .A(n530), .Z(n572) );
  B4I U251 ( .A(n531), .Z(n574) );
  B2I U252 ( .A(data_scrambled[1]), .Z1(n521), .Z2(n533) );
  EN U253 ( .A(n671), .B(n[144]), .Z(data_scrambled[1]) );
  B2I U254 ( .A(n699), .Z1(data_scrambled[4]), .Z2(n532) );
  B2I U255 ( .A(n654), .Z1(), .Z2(n481) );
  IVP U256 ( .A(reset), .Z(n701) );
  B2I U257 ( .A(n661), .Z1(), .Z2(n656) );
  B2I U258 ( .A(n504), .Z1(), .Z2(n659) );
  IVDA U259 ( .A(U4_DATA2_10), .Y(n512), .Z(data_scrambled[16]) );
  EOP U260 ( .A(n684), .B(data_66b_tpg[20]), .Z(n696) );
  IVP U261 ( .A(n696), .Z(data_scrambled[20]) );
  IVDA U262 ( .A(U4_DATA2_0), .Y(n509), .Z(data_scrambled[6]) );
  ENP U263 ( .A(n663), .B(n[149]), .Z(U4_DATA2_0) );
  IVDA U264 ( .A(U4_DATA2_12), .Y(n511), .Z(data_scrambled[18]) );
  ENP U265 ( .A(n667), .B(n497), .Z(U4_DATA2_12) );
  IVDA U266 ( .A(U4_DATA2_5), .Y(n510), .Z(data_scrambled[11]) );
  ENP U267 ( .A(n678), .B(n495), .Z(U4_DATA2_5) );
  ENP U268 ( .A(n681), .B(n[157]), .Z(U4_DATA2_8) );
  IVP U269 ( .A(n490), .Z(n491) );
  IVP U270 ( .A(n492), .Z(n493) );
  IVP U271 ( .A(n494), .Z(n495) );
  IVP U272 ( .A(n496), .Z(n497) );
  IVP U273 ( .A(n498), .Z(n499) );
  EN U274 ( .A(n[144]), .B(n605), .Z(n684) );
  B2I U275 ( .A(n662), .Z1(), .Z2(n500) );
  B2IP U276 ( .A(n662), .Z1(), .Z2(n501) );
  B2IP U277 ( .A(n662), .Z1(), .Z2(n502) );
  B2IP U278 ( .A(n662), .Z1(), .Z2(n503) );
  B5IP U279 ( .A(reset), .Z(n662) );
  B2I U280 ( .A(n500), .Z1(), .Z2(assertion_shengyushen) );
  AN2 U281 ( .A(n577), .B(n578), .Z(n576) );
  AN2 U282 ( .A(n585), .B(n586), .Z(n584) );
  AN2 U283 ( .A(n581), .B(n582), .Z(n580) );
  AN2 U284 ( .A(n589), .B(n590), .Z(n588) );
  IVAP U285 ( .A(n533), .Z(n685) );
  EO U286 ( .A(n593), .B(data_66b_tpg[40]), .Z(data_scrambled[40]) );
  EO U287 ( .A(n525), .B(data_66b_tpg[55]), .Z(data_scrambled[55]) );
  EO U288 ( .A(n518), .B(data_66b_tpg[62]), .Z(data_scrambled[62]) );
  ND2 U289 ( .A(n549), .B(n550), .Z(n518) );
  OR2 U290 ( .A(data_scrambled[20]), .B(n521), .Z(n642) );
  EO U291 ( .A(n596), .B(data_66b_tpg[60]), .Z(data_scrambled[60]) );
  IV U292 ( .A(n616), .Z(n522) );
  ND2 U293 ( .A(data_scrambled[6]), .B(n508), .Z(n523) );
  ND2 U294 ( .A(data_scrambled[11]), .B(n505), .Z(n524) );
  ND2 U295 ( .A(data_scrambled[16]), .B(n507), .Z(n526) );
  ND2 U296 ( .A(n512), .B(n483), .Z(n527) );
  ND2 U297 ( .A(n526), .B(n527), .Z(n525) );
  ND2 U298 ( .A(data_scrambled[18]), .B(n506), .Z(n528) );
  B2IP U299 ( .A(n569), .Z1(n516), .Z2(n529) );
  B2IP U300 ( .A(n571), .Z1(n519), .Z2(n530) );
  B2IP U301 ( .A(n573), .Z1(n517), .Z2(n531) );
  AN2P U302 ( .A(n641), .B(n642), .Z(n640) );
  B2IP U303 ( .A(data_scrambled[0]), .Z1(n480), .Z2(n534) );
  B2IP U304 ( .A(data_scrambled[3]), .Z1(), .Z2(n535) );
  B2IP U305 ( .A(n700), .Z1(), .Z2(data_scrambled[2]) );
  B2IP U306 ( .A(n698), .Z1(), .Z2(data_scrambled[5]) );
  B2I U307 ( .A(n552), .Z1(n473), .Z2(n541) );
  B2I U308 ( .A(n553), .Z1(n475), .Z2(n542) );
  B2I U309 ( .A(n554), .Z1(n477), .Z2(n543) );
  B2I U310 ( .A(n555), .Z1(n469), .Z2(n544) );
  EO1P U311 ( .A(data_scrambled[5]), .B(n471), .C(n470), .D(data_scrambled[5]), 
        .Z(n676) );
  ND2 U312 ( .A(n546), .B(n534), .Z(n545) );
  IV U313 ( .A(data_scrambled[19]), .Z(n546) );
  ND2 U314 ( .A(data_scrambled[22]), .B(n689), .Z(n547) );
  IV U315 ( .A(data_scrambled[22]), .Z(n548) );
  ND2 U316 ( .A(data_scrambled[23]), .B(n532), .Z(n549) );
  ND2 U317 ( .A(n551), .B(data_scrambled[4]), .Z(n550) );
  IV U318 ( .A(data_scrambled[23]), .Z(n551) );
  ENP U319 ( .A(n664), .B(n572), .Z(data_scrambled[7]) );
  ENP U320 ( .A(n[131]), .B(data_66b_tpg[7]), .Z(n664) );
  IV U321 ( .A(n616), .Z(data_scrambled[9]) );
  IVP U322 ( .A(U4_DATA2_3), .Z(n616) );
  ENP U323 ( .A(n680), .B(n570), .Z(data_scrambled[13]) );
  ENP U324 ( .A(n[137]), .B(data_66b_tpg[13]), .Z(n680) );
  ENP U325 ( .A(n679), .B(n574), .Z(data_scrambled[12]) );
  ENP U326 ( .A(n[136]), .B(data_66b_tpg[12]), .Z(n679) );
  ENP U327 ( .A(n[124]), .B(data_66b_tpg[0]), .Z(n670) );
  ENP U328 ( .A(n[127]), .B(data_66b_tpg[3]), .Z(n673) );
  ENP U329 ( .A(n[128]), .B(data_66b_tpg[4]), .Z(n674) );
  ND2 U330 ( .A(n470), .B(n[149]), .Z(n577) );
  ND2 U331 ( .A(n609), .B(n579), .Z(n578) );
  ND2 U332 ( .A(n472), .B(n[151]), .Z(n581) );
  ND2 U333 ( .A(n541), .B(n583), .Z(n582) );
  ND2 U334 ( .A(n474), .B(n[153]), .Z(n585) );
  ND2 U335 ( .A(n542), .B(n587), .Z(n586) );
  ND2 U336 ( .A(n476), .B(n[157]), .Z(n589) );
  ND2 U337 ( .A(n543), .B(n591), .Z(n590) );
  ND2 U338 ( .A(n487), .B(n534), .Z(n592) );
  ND2 U339 ( .A(n608), .B(n685), .Z(n594) );
  ND2 U340 ( .A(n488), .B(n533), .Z(n595) );
  ND2 U341 ( .A(n594), .B(n595), .Z(n593) );
  ND2 U342 ( .A(data_scrambled[21]), .B(n687), .Z(n597) );
  ND2 U343 ( .A(n599), .B(data_scrambled[2]), .Z(n598) );
  IV U344 ( .A(data_scrambled[21]), .Z(n599) );
  ND2 U345 ( .A(n597), .B(n598), .Z(n596) );
  B2I U346 ( .A(n[167]), .Z1(), .Z2(n660) );
  ENP U347 ( .A(n[143]), .B(n670), .Z(data_scrambled[0]) );
  ENP U348 ( .A(n[146]), .B(n673), .Z(data_scrambled[3]) );
  ENP U349 ( .A(n672), .B(n[145]), .Z(n700) );
  B2I U350 ( .A(U4_DATA2_11), .Z1(), .Z2(data_scrambled[17]) );
  EOP U351 ( .A(n690), .B(data_66b_tpg[23]), .Z(n693) );
  IVP U352 ( .A(n693), .Z(data_scrambled[23]) );
  ENP U353 ( .A(n665), .B(n491), .Z(U4_DATA2_10) );
  B2IP U354 ( .A(n500), .Z1(n657), .Z2(n504) );
  ND2 U355 ( .A(data_scrambled[7]), .B(n473), .Z(n614) );
  ND2 U356 ( .A(n522), .B(n475), .Z(n615) );
  ENP U357 ( .A(n669), .B(n493), .Z(U4_DATA2_3) );
  ND2 U358 ( .A(n[166]), .B(n689), .Z(n617) );
  ND2 U359 ( .A(n507), .B(n[160]), .Z(n620) );
  ND2 U360 ( .A(n483), .B(n622), .Z(n621) );
  ND2 U361 ( .A(n620), .B(n621), .Z(n619) );
  ND2 U362 ( .A(n[162]), .B(n506), .Z(n624) );
  ND2 U363 ( .A(n626), .B(n485), .Z(n625) );
  ND2 U364 ( .A(n624), .B(n625), .Z(n623) );
  ND2 U365 ( .A(n468), .B(n516), .Z(n628) );
  ND2 U366 ( .A(n544), .B(n529), .Z(n629) );
  ND2 U367 ( .A(n628), .B(n629), .Z(n627) );
  ND2 U368 ( .A(n508), .B(n519), .Z(n631) );
  ND2 U369 ( .A(n486), .B(n530), .Z(n632) );
  ND2 U370 ( .A(n631), .B(n632), .Z(n630) );
  ND2 U371 ( .A(n[165]), .B(n687), .Z(n633) );
  ND2 U372 ( .A(n505), .B(n517), .Z(n636) );
  ND2 U373 ( .A(n484), .B(n531), .Z(n637) );
  ND2 U374 ( .A(n636), .B(n637), .Z(n635) );
  ND2 U375 ( .A(data_scrambled[13]), .B(n477), .Z(n638) );
  ND2 U376 ( .A(data_scrambled[12]), .B(n469), .Z(n639) );
  ND2 U377 ( .A(data_scrambled[20]), .B(n685), .Z(n641) );
  B2I U378 ( .A(U4_DATA2_9), .Z1(), .Z2(data_scrambled[15]) );
  EOP U379 ( .A(n686), .B(data_66b_tpg[21]), .Z(n695) );
  IVP U380 ( .A(n695), .Z(data_scrambled[21]) );
  B2I U381 ( .A(U4_DATA2_8), .Z1(), .Z2(data_scrambled[14]) );
  B2I U382 ( .A(U4_DATA2_2), .Z1(), .Z2(data_scrambled[8]) );
  EOP U383 ( .A(n688), .B(data_66b_tpg[22]), .Z(n694) );
  IVP U384 ( .A(n694), .Z(data_scrambled[22]) );
  B2I U385 ( .A(U4_DATA2_4), .Z1(), .Z2(data_scrambled[10]) );
  EOP U386 ( .A(n683), .B(data_66b_tpg[19]), .Z(n697) );
  IVP U387 ( .A(n697), .Z(data_scrambled[19]) );
  ENP U388 ( .A(n675), .B(n[148]), .Z(n698) );
  IVP U389 ( .A(n657), .Z(n661) );
  EN U390 ( .A(n[130]), .B(data_66b_tpg[6]), .Z(n663) );
  EN U391 ( .A(n[140]), .B(data_66b_tpg[16]), .Z(n665) );
  EN U392 ( .A(n[141]), .B(data_66b_tpg[17]), .Z(n666) );
  EN U393 ( .A(n666), .B(n[160]), .Z(U4_DATA2_11) );
  EN U394 ( .A(n[142]), .B(data_66b_tpg[18]), .Z(n667) );
  EN U395 ( .A(n576), .B(data_66b_tpg[25]), .Z(data_scrambled[25]) );
  EN U396 ( .A(data_66b_tpg[8]), .B(n[132]), .Z(n668) );
  EN U397 ( .A(n668), .B(n[151]), .Z(U4_DATA2_2) );
  EN U398 ( .A(n580), .B(data_66b_tpg[27]), .Z(data_scrambled[27]) );
  EN U399 ( .A(n584), .B(data_66b_tpg[29]), .Z(data_scrambled[29]) );
  EN U400 ( .A(n588), .B(data_66b_tpg[33]), .Z(data_scrambled[33]) );
  EN U401 ( .A(n[129]), .B(data_66b_tpg[5]), .Z(n675) );
  EN U402 ( .A(n676), .B(data_66b_tpg[44]), .Z(data_scrambled[44]) );
  EN U403 ( .A(n[134]), .B(data_66b_tpg[10]), .Z(n677) );
  EN U404 ( .A(n677), .B(n[153]), .Z(U4_DATA2_4) );
  EN U405 ( .A(n[135]), .B(data_66b_tpg[11]), .Z(n678) );
  EN U406 ( .A(n[138]), .B(data_66b_tpg[14]), .Z(n681) );
  EN U407 ( .A(n[139]), .B(data_66b_tpg[15]), .Z(n682) );
  EN U408 ( .A(n682), .B(n499), .Z(U4_DATA2_9) );
  EN U409 ( .A(n[162]), .B(n[143]), .Z(n683) );
  EN U410 ( .A(n[145]), .B(n608), .Z(n686) );
  EN U411 ( .A(n[165]), .B(n[146]), .Z(n688) );
  EN U412 ( .A(n[166]), .B(n[147]), .Z(n690) );
  EN U413 ( .A(n[148]), .B(n[167]), .Z(n691) );
endmodule

