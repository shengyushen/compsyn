
module XFIPCS_64B66B_ENC ( CLK, RESET, DATA_VALID, ENCODER_DATA_IN, 
        ENCODER_CONTROL_IN, TEST_PAT_SEED_A, TEST_PAT_SEED_B, TEST_MODE, 
        DATA_PAT_SEL, ENCODER_DATA_OUT, assertion_shengyushen );
  input [63:0] ENCODER_DATA_IN;
  input [7:0] ENCODER_CONTROL_IN;
  input [57:0] TEST_PAT_SEED_A;
  input [57:0] TEST_PAT_SEED_B;
  output [65:0] ENCODER_DATA_OUT;
  input CLK, RESET, DATA_VALID, TEST_MODE, DATA_PAT_SEL;
  output assertion_shengyushen;
  wire   n3, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n278, n279, n281, n283, n284, n286, n287, n289, n290,
         n295, n296, n297, n301, n305, n306, n308, n309, n310, n314, n316,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n919, n920, n921, n922, n923,
         n924, n925, n926, n931, n932, n933, n934, n935, n936, n937, n938,
         n940, n941, n942, n943, n944, n945, n946, n947, n949, n950, n951,
         n952, n953, n954, n955, n956, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n1046, n1057, n1062, n1237, n1296,
         n1297, n1363, n1364, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1781, n1783, n1785, n1787, n1789,
         n1791, n1793, n1795, n1797, n1799, n1801, n1803, n1805, n1807, n1809,
         n1811, n1813, n1815, n1817, n1819, n1821, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1970, n1971,
         U3_n725, U34_Z_0, U34_Z_1, U34_Z_2, U34_CONTROL2, U34_CONTROL1,
         U34_DATA1_0, U34_DATA1_1, U34_DATA1_2, U33_Z_0, U33_Z_1, U33_Z_2,
         U33_Z_3, U33_CONTROL5, U33_DATA1_0, U33_DATA1_1, U33_DATA1_2,
         U33_DATA1_3, U32_Z_0, U32_CONTROL1, U32_DATA1_0, U31_Z_0, U31_Z_1,
         U31_Z_2, U31_Z_3, U31_DATA1_0, U31_DATA1_1, U31_DATA1_2, U31_DATA1_3,
         U30_Z_0, U30_Z_1, U30_DATA1_0, U30_DATA1_1, U29_Z_0, U29_Z_1,
         U29_CONTROL1, U29_DATA1_0, U29_DATA1_1, U28_Z_0, U28_Z_1, U28_Z_2,
         U28_CONTROL4, U28_DATA1_0, U28_DATA1_1, U28_DATA1_2, U27_Z_0, U27_Z_1,
         U27_DATA1_0, U27_DATA1_1, U26_Z_0, U26_Z_1, U26_Z_2, U26_DATA1_0,
         U26_DATA1_1, U26_DATA1_2, U25_Z_0, U25_Z_1, U25_CONTROL5,
         U25_CONTROL2, U25_DATA1_0, U25_DATA1_1, U24_Z_0, U24_Z_1, U24_DATA1_0,
         U24_DATA1_1, U23_Z_0, U23_DATA1_0, U20_Z_0, U20_Z_1, U20_Z_2,
         U20_DATA1_0, U20_DATA1_1, U20_DATA1_2, U19_Z_0, U19_CONTROL4,
         U19_CONTROL2, U19_DATA1_0, U18_Z_0, U18_Z_1, U18_DATA1_0, U18_DATA1_1,
         U17_Z_0, U17_Z_1, U17_Z_2, U17_Z_3, U17_Z_4, U17_DATA1_0, U17_DATA1_1,
         U17_DATA1_2, U17_DATA1_3, U17_DATA1_4, U16_Z_0, U16_Z_1, U16_DATA1_0,
         U16_DATA1_1, U15_Z_0, U15_Z_1, U15_Z_2, U15_Z_3, U15_Z_4, U15_Z_5,
         U15_DATA1_0, U15_DATA1_1, U15_DATA1_2, U15_DATA1_3, U15_DATA1_4,
         U15_DATA1_5, U14_Z_0, U14_DATA1_0, U13_Z_0, U13_Z_1, U13_Z_2, U13_Z_3,
         U13_Z_4, U13_Z_5, U13_Z_6, U13_DATA1_0, U13_DATA1_1, U13_DATA1_2,
         U13_DATA1_3, U13_DATA1_4, U13_DATA1_5, U13_DATA1_6, U10_DATA2_0,
         U10_DATA2_1, U10_DATA2_2, U10_DATA2_3, U10_DATA2_4, U10_DATA2_5,
         U10_DATA2_6, U10_DATA2_7, U7_DATA6_0, U7_DATA6_1, U7_DATA6_2,
         U7_DATA6_3, U7_DATA6_4, U7_DATA6_5, U7_DATA6_6, U7_DATA6_7,
         U7_DATA6_8, U7_DATA6_9, U7_DATA6_10, U7_DATA6_11, U7_DATA6_12,
         U7_DATA6_13, U7_DATA6_14, U7_DATA6_15, U7_DATA6_16, U7_DATA6_17,
         U7_DATA6_18, U7_DATA6_19, U7_DATA6_20, U7_DATA6_21, U7_DATA6_22,
         U7_DATA6_23, U7_DATA6_24, U7_DATA6_25, U7_DATA6_26, U7_DATA6_27,
         U7_DATA6_28, U7_DATA6_29, U7_DATA6_30, U7_DATA6_31, U7_DATA6_32,
         U7_DATA6_33, U7_DATA6_34, U7_DATA6_35, U7_DATA6_36, U7_DATA6_37,
         U7_DATA6_38, U7_DATA6_39, U7_DATA6_40, U7_DATA6_41, U7_DATA6_42,
         U7_DATA6_43, U7_DATA6_44, U7_DATA6_45, U7_DATA6_46, U7_DATA6_47,
         U7_DATA6_48, U7_DATA6_49, U7_DATA6_50, U7_DATA6_51, U7_DATA6_52,
         U7_DATA6_53, U7_DATA6_54, U7_DATA6_55, U7_DATA6_56, U7_DATA6_57,
         U7_DATA4_0, U7_DATA4_1, U7_DATA4_2, U7_DATA4_3, U7_DATA4_4,
         U7_DATA4_5, U7_DATA4_6, U7_DATA4_7, U7_DATA4_8, U7_DATA4_9,
         U7_DATA4_10, U7_DATA4_11, U7_DATA4_12, U7_DATA4_13, U7_DATA4_14,
         U7_DATA4_15, U7_DATA4_16, U7_DATA4_17, U7_DATA4_18, U7_DATA4_19,
         U7_DATA4_20, U7_DATA4_21, U7_DATA4_22, U7_DATA4_23, U7_DATA4_24,
         U7_DATA4_25, U7_DATA4_26, U7_DATA4_27, U7_DATA4_28, U7_DATA4_29,
         U7_DATA4_30, U7_DATA4_31, U7_DATA4_32, U7_DATA4_33, U7_DATA4_34,
         U7_DATA4_35, U7_DATA4_36, U7_DATA4_37, U7_DATA4_38, U7_DATA4_39,
         U7_DATA4_40, U7_DATA4_41, U7_DATA4_42, U7_DATA4_43, U7_DATA4_44,
         U7_DATA4_45, U7_DATA4_46, U7_DATA4_47, U7_DATA4_48, U7_DATA4_49,
         U7_DATA4_50, U7_DATA4_51, U7_DATA4_52, U7_DATA4_53, U7_DATA4_54,
         U7_DATA4_55, U7_DATA4_56, U7_DATA4_57, U7_DATA1_0, U7_DATA1_1,
         U7_DATA1_2, U7_DATA1_3, U7_DATA1_4, U7_DATA1_5, U7_DATA1_6,
         U7_DATA1_7, U7_DATA1_8, U7_DATA1_9, U7_DATA1_10, U7_DATA1_11,
         U7_DATA1_12, U7_DATA1_13, U7_DATA1_14, U7_DATA1_15, U7_DATA1_16,
         U7_DATA1_17, U7_DATA1_18, U7_DATA1_19, U7_DATA1_20, U7_DATA1_21,
         U7_DATA1_22, U7_DATA1_23, U7_DATA1_24, U7_DATA1_25, U7_DATA1_26,
         U7_DATA1_27, U7_DATA1_28, U7_DATA1_29, U7_DATA1_30, U7_DATA1_31,
         U7_DATA1_32, U7_DATA1_33, U7_DATA1_34, U7_DATA1_35, U7_DATA1_36,
         U7_DATA1_37, U7_DATA1_38, U7_DATA1_39, U7_DATA1_40, U7_DATA1_41,
         U7_DATA1_42, U7_DATA1_43, U7_DATA1_44, U7_DATA1_45, U7_DATA1_46,
         U7_DATA1_47, U7_DATA1_48, U7_DATA1_49, U7_DATA1_50, U7_DATA1_51,
         U7_DATA1_52, U7_DATA1_53, U7_DATA1_54, U7_DATA1_55, U7_DATA1_56,
         U7_DATA1_57, U6_Z_0, U6_Z_1, U6_Z_2, U6_Z_3, U6_Z_4, U6_Z_5, U6_Z_6,
         U6_Z_7, U6_Z_8, U5_Z_0, U5_Z_1, U5_Z_2, U5_Z_3, U5_Z_4, U5_Z_5,
         U5_Z_6, U5_Z_7, U5_Z_8, U5_Z_9, U5_Z_10, U5_Z_11, U5_Z_12, U5_Z_13,
         U5_Z_14, U5_Z_15, U5_Z_16, U5_Z_17, U5_Z_18, U5_Z_19, U5_Z_20,
         U5_Z_21, U5_Z_22, U5_Z_23, U5_Z_24, U5_Z_25, U5_Z_26, U5_Z_27,
         U5_Z_28, U5_Z_29, U5_Z_30, U5_Z_31, U5_Z_32, U5_Z_33, U5_Z_34,
         U5_Z_35, U5_Z_36, U5_Z_37, U5_Z_38, U5_Z_39, U5_Z_40, U5_Z_41,
         U5_Z_42, U5_Z_43, U5_Z_44, U5_Z_45, U5_Z_46, U5_Z_47, U5_Z_48,
         U5_Z_49, U5_Z_50, U5_Z_51, U5_Z_52, U5_Z_53, U5_Z_54, U5_Z_55,
         U5_Z_56, U5_Z_57, U4_DATA1_0, U4_DATA1_1, U4_DATA1_2, U4_DATA1_3,
         U4_DATA1_4, U4_DATA1_5, U4_DATA1_6, U4_DATA1_7, U4_DATA1_8, n2412,
         n2460, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2491, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2661, n3749, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760;
  wire   [1757:1743] n;

  AN2 C6836 ( .A(n969), .B(n968), .Z(n8) );
  AN2 C6835 ( .A(n8), .B(n967), .Z(n7) );
  AN2 C6834 ( .A(n7), .B(DATA_VALID), .Z(assertion_shengyushen) );
  OR2 C6833 ( .A(n[1757]), .B(n[1756]), .Z(n22) );
  OR2 C6832 ( .A(n22), .B(n[1755]), .Z(n21) );
  OR2 C6831 ( .A(n21), .B(n[1754]), .Z(n20) );
  OR2 C6830 ( .A(n20), .B(n[1753]), .Z(n19) );
  OR2 C6829 ( .A(n19), .B(n[1752]), .Z(n18) );
  OR2 C6828 ( .A(n18), .B(n[1751]), .Z(n17) );
  OR2 C6827 ( .A(n17), .B(n[1750]), .Z(n16) );
  OR2 C6826 ( .A(n16), .B(n[1749]), .Z(n15) );
  OR2 C6825 ( .A(n15), .B(n[1748]), .Z(n14) );
  OR2 C6824 ( .A(n14), .B(n[1747]), .Z(n13) );
  OR2 C6823 ( .A(n13), .B(n[1746]), .Z(n12) );
  OR2 C6822 ( .A(n12), .B(n[1745]), .Z(n11) );
  OR2 C6821 ( .A(n11), .B(n[1744]), .Z(n10) );
  OR2 C6820 ( .A(n10), .B(n[1743]), .Z(n9) );
  OR2 C6819 ( .A(n9), .B(n959), .Z(n969) );
  IV I_346 ( .A(DATA_VALID), .Z(n1046) );
  OR2 C6807 ( .A(RESET), .B(n2491), .Z(n1057) );
  IV I_344 ( .A(TEST_PAT_SEED_B[0]), .Z(U7_DATA6_0) );
  IV I_343 ( .A(TEST_PAT_SEED_B[1]), .Z(U7_DATA6_1) );
  IV I_342 ( .A(TEST_PAT_SEED_B[2]), .Z(U7_DATA6_2) );
  IV I_341 ( .A(TEST_PAT_SEED_B[3]), .Z(U7_DATA6_3) );
  IV I_340 ( .A(TEST_PAT_SEED_B[4]), .Z(U7_DATA6_4) );
  IV I_339 ( .A(TEST_PAT_SEED_B[5]), .Z(U7_DATA6_5) );
  IV I_338 ( .A(TEST_PAT_SEED_B[6]), .Z(U7_DATA6_6) );
  IV I_337 ( .A(TEST_PAT_SEED_B[7]), .Z(U7_DATA6_7) );
  IV I_336 ( .A(TEST_PAT_SEED_B[8]), .Z(U7_DATA6_8) );
  IV I_335 ( .A(TEST_PAT_SEED_B[9]), .Z(U7_DATA6_9) );
  IV I_334 ( .A(TEST_PAT_SEED_B[10]), .Z(U7_DATA6_10) );
  IV I_333 ( .A(TEST_PAT_SEED_B[11]), .Z(U7_DATA6_11) );
  IV I_332 ( .A(TEST_PAT_SEED_B[12]), .Z(U7_DATA6_12) );
  IV I_331 ( .A(TEST_PAT_SEED_B[13]), .Z(U7_DATA6_13) );
  IV I_330 ( .A(TEST_PAT_SEED_B[14]), .Z(U7_DATA6_14) );
  IV I_329 ( .A(TEST_PAT_SEED_B[15]), .Z(U7_DATA6_15) );
  IV I_328 ( .A(TEST_PAT_SEED_B[16]), .Z(U7_DATA6_16) );
  IV I_327 ( .A(TEST_PAT_SEED_B[17]), .Z(U7_DATA6_17) );
  IV I_326 ( .A(TEST_PAT_SEED_B[18]), .Z(U7_DATA6_18) );
  IV I_325 ( .A(TEST_PAT_SEED_B[19]), .Z(U7_DATA6_19) );
  IV I_324 ( .A(TEST_PAT_SEED_B[20]), .Z(U7_DATA6_20) );
  IV I_323 ( .A(TEST_PAT_SEED_B[21]), .Z(U7_DATA6_21) );
  IV I_322 ( .A(TEST_PAT_SEED_B[22]), .Z(U7_DATA6_22) );
  IV I_321 ( .A(TEST_PAT_SEED_B[23]), .Z(U7_DATA6_23) );
  IV I_320 ( .A(TEST_PAT_SEED_B[24]), .Z(U7_DATA6_24) );
  IV I_319 ( .A(TEST_PAT_SEED_B[25]), .Z(U7_DATA6_25) );
  IV I_318 ( .A(TEST_PAT_SEED_B[26]), .Z(U7_DATA6_26) );
  IV I_317 ( .A(TEST_PAT_SEED_B[27]), .Z(U7_DATA6_27) );
  IV I_316 ( .A(TEST_PAT_SEED_B[28]), .Z(U7_DATA6_28) );
  IV I_315 ( .A(TEST_PAT_SEED_B[29]), .Z(U7_DATA6_29) );
  IV I_314 ( .A(TEST_PAT_SEED_B[30]), .Z(U7_DATA6_30) );
  IV I_313 ( .A(TEST_PAT_SEED_B[31]), .Z(U7_DATA6_31) );
  IV I_312 ( .A(TEST_PAT_SEED_B[32]), .Z(U7_DATA6_32) );
  IV I_311 ( .A(TEST_PAT_SEED_B[33]), .Z(U7_DATA6_33) );
  IV I_310 ( .A(TEST_PAT_SEED_B[34]), .Z(U7_DATA6_34) );
  IV I_309 ( .A(TEST_PAT_SEED_B[35]), .Z(U7_DATA6_35) );
  IV I_308 ( .A(TEST_PAT_SEED_B[36]), .Z(U7_DATA6_36) );
  IV I_307 ( .A(TEST_PAT_SEED_B[37]), .Z(U7_DATA6_37) );
  IV I_306 ( .A(TEST_PAT_SEED_B[38]), .Z(U7_DATA6_38) );
  IV I_305 ( .A(TEST_PAT_SEED_B[39]), .Z(U7_DATA6_39) );
  IV I_304 ( .A(TEST_PAT_SEED_B[40]), .Z(U7_DATA6_40) );
  IV I_303 ( .A(TEST_PAT_SEED_B[41]), .Z(U7_DATA6_41) );
  IV I_302 ( .A(TEST_PAT_SEED_B[42]), .Z(U7_DATA6_42) );
  IV I_301 ( .A(TEST_PAT_SEED_B[43]), .Z(U7_DATA6_43) );
  IV I_300 ( .A(TEST_PAT_SEED_B[44]), .Z(U7_DATA6_44) );
  IV I_299 ( .A(TEST_PAT_SEED_B[45]), .Z(U7_DATA6_45) );
  IV I_298 ( .A(TEST_PAT_SEED_B[46]), .Z(U7_DATA6_46) );
  IV I_297 ( .A(TEST_PAT_SEED_B[47]), .Z(U7_DATA6_47) );
  IV I_296 ( .A(TEST_PAT_SEED_B[48]), .Z(U7_DATA6_48) );
  IV I_295 ( .A(TEST_PAT_SEED_B[49]), .Z(U7_DATA6_49) );
  IV I_294 ( .A(TEST_PAT_SEED_B[50]), .Z(U7_DATA6_50) );
  IV I_293 ( .A(TEST_PAT_SEED_B[51]), .Z(U7_DATA6_51) );
  IV I_292 ( .A(TEST_PAT_SEED_B[52]), .Z(U7_DATA6_52) );
  IV I_291 ( .A(TEST_PAT_SEED_B[53]), .Z(U7_DATA6_53) );
  IV I_290 ( .A(TEST_PAT_SEED_B[54]), .Z(U7_DATA6_54) );
  IV I_289 ( .A(TEST_PAT_SEED_B[55]), .Z(U7_DATA6_55) );
  IV I_288 ( .A(TEST_PAT_SEED_B[56]), .Z(U7_DATA6_56) );
  IV I_287 ( .A(TEST_PAT_SEED_B[57]), .Z(U7_DATA6_57) );
  IV I_286 ( .A(TEST_PAT_SEED_A[0]), .Z(U7_DATA4_0) );
  IV I_285 ( .A(TEST_PAT_SEED_A[1]), .Z(U7_DATA4_1) );
  IV I_284 ( .A(TEST_PAT_SEED_A[2]), .Z(U7_DATA4_2) );
  IV I_283 ( .A(TEST_PAT_SEED_A[3]), .Z(U7_DATA4_3) );
  IV I_282 ( .A(TEST_PAT_SEED_A[4]), .Z(U7_DATA4_4) );
  IV I_281 ( .A(TEST_PAT_SEED_A[5]), .Z(U7_DATA4_5) );
  IV I_280 ( .A(TEST_PAT_SEED_A[6]), .Z(U7_DATA4_6) );
  IV I_279 ( .A(TEST_PAT_SEED_A[7]), .Z(U7_DATA4_7) );
  IV I_278 ( .A(TEST_PAT_SEED_A[8]), .Z(U7_DATA4_8) );
  IV I_277 ( .A(TEST_PAT_SEED_A[9]), .Z(U7_DATA4_9) );
  IV I_276 ( .A(TEST_PAT_SEED_A[10]), .Z(U7_DATA4_10) );
  IV I_275 ( .A(TEST_PAT_SEED_A[11]), .Z(U7_DATA4_11) );
  IV I_274 ( .A(TEST_PAT_SEED_A[12]), .Z(U7_DATA4_12) );
  IV I_273 ( .A(TEST_PAT_SEED_A[13]), .Z(U7_DATA4_13) );
  IV I_272 ( .A(TEST_PAT_SEED_A[14]), .Z(U7_DATA4_14) );
  IV I_271 ( .A(TEST_PAT_SEED_A[15]), .Z(U7_DATA4_15) );
  IV I_270 ( .A(TEST_PAT_SEED_A[16]), .Z(U7_DATA4_16) );
  IV I_269 ( .A(TEST_PAT_SEED_A[17]), .Z(U7_DATA4_17) );
  IV I_268 ( .A(TEST_PAT_SEED_A[18]), .Z(U7_DATA4_18) );
  IV I_267 ( .A(TEST_PAT_SEED_A[19]), .Z(U7_DATA4_19) );
  IV I_266 ( .A(TEST_PAT_SEED_A[20]), .Z(U7_DATA4_20) );
  IV I_265 ( .A(TEST_PAT_SEED_A[21]), .Z(U7_DATA4_21) );
  IV I_264 ( .A(TEST_PAT_SEED_A[22]), .Z(U7_DATA4_22) );
  IV I_263 ( .A(TEST_PAT_SEED_A[23]), .Z(U7_DATA4_23) );
  IV I_262 ( .A(TEST_PAT_SEED_A[24]), .Z(U7_DATA4_24) );
  IV I_261 ( .A(TEST_PAT_SEED_A[25]), .Z(U7_DATA4_25) );
  IV I_260 ( .A(TEST_PAT_SEED_A[26]), .Z(U7_DATA4_26) );
  IV I_259 ( .A(TEST_PAT_SEED_A[27]), .Z(U7_DATA4_27) );
  IV I_258 ( .A(TEST_PAT_SEED_A[28]), .Z(U7_DATA4_28) );
  IV I_257 ( .A(TEST_PAT_SEED_A[29]), .Z(U7_DATA4_29) );
  IV I_256 ( .A(TEST_PAT_SEED_A[30]), .Z(U7_DATA4_30) );
  IV I_255 ( .A(TEST_PAT_SEED_A[31]), .Z(U7_DATA4_31) );
  IV I_254 ( .A(TEST_PAT_SEED_A[32]), .Z(U7_DATA4_32) );
  IV I_253 ( .A(TEST_PAT_SEED_A[33]), .Z(U7_DATA4_33) );
  IV I_252 ( .A(TEST_PAT_SEED_A[34]), .Z(U7_DATA4_34) );
  IV I_251 ( .A(TEST_PAT_SEED_A[35]), .Z(U7_DATA4_35) );
  IV I_250 ( .A(TEST_PAT_SEED_A[36]), .Z(U7_DATA4_36) );
  IV I_249 ( .A(TEST_PAT_SEED_A[37]), .Z(U7_DATA4_37) );
  IV I_248 ( .A(TEST_PAT_SEED_A[38]), .Z(U7_DATA4_38) );
  IV I_247 ( .A(TEST_PAT_SEED_A[39]), .Z(U7_DATA4_39) );
  IV I_246 ( .A(TEST_PAT_SEED_A[40]), .Z(U7_DATA4_40) );
  IV I_245 ( .A(TEST_PAT_SEED_A[41]), .Z(U7_DATA4_41) );
  IV I_244 ( .A(TEST_PAT_SEED_A[42]), .Z(U7_DATA4_42) );
  IV I_243 ( .A(TEST_PAT_SEED_A[43]), .Z(U7_DATA4_43) );
  IV I_242 ( .A(TEST_PAT_SEED_A[44]), .Z(U7_DATA4_44) );
  IV I_241 ( .A(TEST_PAT_SEED_A[45]), .Z(U7_DATA4_45) );
  IV I_240 ( .A(TEST_PAT_SEED_A[46]), .Z(U7_DATA4_46) );
  IV I_239 ( .A(TEST_PAT_SEED_A[47]), .Z(U7_DATA4_47) );
  IV I_238 ( .A(TEST_PAT_SEED_A[48]), .Z(U7_DATA4_48) );
  IV I_237 ( .A(TEST_PAT_SEED_A[49]), .Z(U7_DATA4_49) );
  IV I_236 ( .A(TEST_PAT_SEED_A[50]), .Z(U7_DATA4_50) );
  IV I_235 ( .A(TEST_PAT_SEED_A[51]), .Z(U7_DATA4_51) );
  IV I_234 ( .A(TEST_PAT_SEED_A[52]), .Z(U7_DATA4_52) );
  IV I_233 ( .A(TEST_PAT_SEED_A[53]), .Z(U7_DATA4_53) );
  IV I_232 ( .A(TEST_PAT_SEED_A[54]), .Z(U7_DATA4_54) );
  IV I_231 ( .A(TEST_PAT_SEED_A[55]), .Z(U7_DATA4_55) );
  IV I_230 ( .A(TEST_PAT_SEED_A[56]), .Z(U7_DATA4_56) );
  IV I_229 ( .A(TEST_PAT_SEED_A[57]), .Z(U7_DATA4_57) );
  AN2 C6520 ( .A(n1971), .B(n2460), .Z(n1364) );
  IV I_223 ( .A(n1440), .Z(n1439) );
  IV I_222 ( .A(n[1757]), .Z(n1454) );
  IV I_221 ( .A(n1456), .Z(n1455) );
  IV I_220 ( .A(n[1756]), .Z(n1470) );
  IV I_219 ( .A(n1472), .Z(n1471) );
  IV I_218 ( .A(n[1755]), .Z(n1486) );
  IV I_217 ( .A(n1488), .Z(n1487) );
  IV I_216 ( .A(n[1754]), .Z(n1502) );
  IV I_215 ( .A(n1504), .Z(n1503) );
  IV I_214 ( .A(n[1753]), .Z(n1518) );
  IV I_213 ( .A(n1520), .Z(n1519) );
  IV I_212 ( .A(n[1752]), .Z(n1534) );
  IV I_211 ( .A(n1536), .Z(n1535) );
  IV I_210 ( .A(n[1751]), .Z(n1550) );
  IV I_209 ( .A(n1552), .Z(n1551) );
  IV I_208 ( .A(n[1750]), .Z(n1566) );
  IV I_207 ( .A(n1568), .Z(n1567) );
  IV I_206 ( .A(n[1749]), .Z(n1582) );
  IV I_205 ( .A(n1584), .Z(n1583) );
  IV I_204 ( .A(n[1748]), .Z(n1598) );
  IV I_203 ( .A(n1600), .Z(n1599) );
  IV I_202 ( .A(n[1747]), .Z(n1614) );
  IV I_201 ( .A(n1616), .Z(n1615) );
  IV I_200 ( .A(n[1746]), .Z(n1630) );
  IV I_199 ( .A(n1632), .Z(n1631) );
  IV I_198 ( .A(n[1745]), .Z(n1646) );
  IV I_197 ( .A(n1648), .Z(n1647) );
  IV I_196 ( .A(n[1744]), .Z(n1662) );
  IV I_195 ( .A(n1664), .Z(n1663) );
  IV I_194 ( .A(n[1743]), .Z(n1678) );
  AN2 C6395 ( .A(n1773), .B(n1962), .Z(n87) );
  AN2 C6394 ( .A(n87), .B(n1809), .Z(n1758) );
  AN2 C6393 ( .A(n1773), .B(n1811), .Z(n88) );
  AN2 C6392 ( .A(n88), .B(n1781), .Z(n1759) );
  AN2 C6391 ( .A(n1774), .B(n1813), .Z(n90) );
  AN2 C6390 ( .A(n90), .B(n1783), .Z(n89) );
  AN2 C6389 ( .A(n89), .B(n1781), .Z(n1760) );
  AN2 C6388 ( .A(n1775), .B(n1815), .Z(n93) );
  AN2 C6387 ( .A(n93), .B(n1785), .Z(n92) );
  AN2 C6386 ( .A(n92), .B(n1783), .Z(n91) );
  AN2 C6385 ( .A(n91), .B(n1781), .Z(n1761) );
  AN2 C6384 ( .A(n1776), .B(n1817), .Z(n97) );
  AN2 C6383 ( .A(n97), .B(n1787), .Z(n96) );
  AN2 C6382 ( .A(n96), .B(n1785), .Z(n95) );
  AN2 C6381 ( .A(n95), .B(n1783), .Z(n94) );
  AN2 C6380 ( .A(n94), .B(n1781), .Z(n1762) );
  AN2 C6379 ( .A(n1777), .B(n1819), .Z(n102) );
  AN2 C6378 ( .A(n102), .B(n1789), .Z(n101) );
  AN2 C6377 ( .A(n101), .B(n1787), .Z(n100) );
  AN2 C6376 ( .A(n100), .B(n1785), .Z(n99) );
  AN2 C6375 ( .A(n99), .B(n1783), .Z(n98) );
  AN2 C6374 ( .A(n98), .B(n1781), .Z(n1763) );
  AN2 C6373 ( .A(n1968), .B(n1821), .Z(n108) );
  AN2 C6372 ( .A(n108), .B(n1791), .Z(n107) );
  AN2 C6371 ( .A(n107), .B(n1789), .Z(n106) );
  AN2 C6370 ( .A(n106), .B(n1787), .Z(n105) );
  AN2 C6369 ( .A(n105), .B(n1785), .Z(n104) );
  AN2 C6368 ( .A(n104), .B(n1783), .Z(n103) );
  AN2 C6367 ( .A(n103), .B(n1781), .Z(n1764) );
  AN2 C6366 ( .A(n1823), .B(n1793), .Z(n114) );
  AN2 C6365 ( .A(n114), .B(n1791), .Z(n113) );
  AN2 C6364 ( .A(n113), .B(n1789), .Z(n112) );
  AN2 C6363 ( .A(n112), .B(n1787), .Z(n111) );
  AN2 C6362 ( .A(n111), .B(n1785), .Z(n110) );
  AN2 C6361 ( .A(n110), .B(n1783), .Z(n109) );
  AN2 C6360 ( .A(n109), .B(n1781), .Z(n1765) );
  AN2 C6359 ( .A(n1778), .B(n1787), .Z(n117) );
  AN2 C6358 ( .A(n117), .B(n1785), .Z(n116) );
  AN2 C6357 ( .A(n116), .B(n1783), .Z(n115) );
  AN2 C6356 ( .A(n115), .B(n1781), .Z(n1766) );
  AN2 C6355 ( .A(n1799), .B(n1967), .Z(n123) );
  AN2 C6354 ( .A(n123), .B(n1966), .Z(n122) );
  AN2 C6353 ( .A(n122), .B(n1965), .Z(n121) );
  AN2 C6352 ( .A(n121), .B(n1964), .Z(n120) );
  AN2 C6351 ( .A(n120), .B(n1963), .Z(n119) );
  AN2 C6350 ( .A(n119), .B(n1962), .Z(n118) );
  AN2 C6349 ( .A(n118), .B(n1961), .Z(n1767) );
  AN2 C6348 ( .A(n1778), .B(n1803), .Z(n126) );
  AN2 C6347 ( .A(n126), .B(n1963), .Z(n125) );
  AN2 C6346 ( .A(n125), .B(n1962), .Z(n124) );
  AN2 C6345 ( .A(n124), .B(n1961), .Z(n1768) );
  AN2 C6344 ( .A(n1778), .B(n1797), .Z(n129) );
  AN2 C6343 ( .A(n129), .B(n1963), .Z(n128) );
  AN2 C6342 ( .A(n128), .B(n1962), .Z(n127) );
  AN2 C6341 ( .A(n127), .B(n1961), .Z(n1769) );
  AN2 C6340 ( .A(n1779), .B(n1797), .Z(n132) );
  AN2 C6339 ( .A(n132), .B(n1963), .Z(n131) );
  AN2 C6338 ( .A(n131), .B(n1962), .Z(n130) );
  AN2 C6337 ( .A(n130), .B(n1961), .Z(n1770) );
  AN2 C6336 ( .A(n1779), .B(n1803), .Z(n135) );
  AN2 C6335 ( .A(n135), .B(n1963), .Z(n134) );
  AN2 C6334 ( .A(n134), .B(n1962), .Z(n133) );
  AN2 C6333 ( .A(n133), .B(n1961), .Z(n1771) );
  AN2 C6332 ( .A(n1779), .B(n1787), .Z(n138) );
  AN2 C6331 ( .A(n138), .B(n1785), .Z(n137) );
  AN2 C6330 ( .A(n137), .B(n1783), .Z(n136) );
  AN2 C6329 ( .A(n136), .B(n1781), .Z(n1772) );
  AN2 C6328 ( .A(n1774), .B(n1963), .Z(n1773) );
  AN2 C6327 ( .A(n1775), .B(n1964), .Z(n1774) );
  AN2 C6326 ( .A(n1776), .B(n1965), .Z(n1775) );
  AN2 C6325 ( .A(n1777), .B(n1966), .Z(n1776) );
  AN2 C6324 ( .A(n1968), .B(n1967), .Z(n1777) );
  AN2 C6323 ( .A(n1807), .B(n1967), .Z(n140) );
  AN2 C6322 ( .A(n140), .B(n1966), .Z(n139) );
  AN2 C6321 ( .A(n139), .B(n1965), .Z(n1778) );
  AN2 C6320 ( .A(n1795), .B(n1793), .Z(n142) );
  AN2 C6319 ( .A(n142), .B(n1791), .Z(n141) );
  AN2 C6318 ( .A(n141), .B(n1789), .Z(n1779) );
  OR2 C6316 ( .A(n441), .B(n502), .Z(n149) );
  OR2 C6315 ( .A(n149), .B(n623), .Z(n148) );
  OR2 C6314 ( .A(n148), .B(n564), .Z(n147) );
  OR2 C6313 ( .A(n147), .B(n684), .Z(n146) );
  OR2 C6312 ( .A(n146), .B(n739), .Z(n145) );
  OR2 C6311 ( .A(n145), .B(n802), .Z(n144) );
  OR2 C6310 ( .A(n144), .B(n903), .Z(n143) );
  AN2 C6309 ( .A(ENCODER_CONTROL_IN[7]), .B(n143), .Z(n1781) );
  OR2 C6307 ( .A(n426), .B(n486), .Z(n156) );
  OR2 C6306 ( .A(n156), .B(n608), .Z(n155) );
  OR2 C6305 ( .A(n155), .B(n549), .Z(n154) );
  OR2 C6304 ( .A(n154), .B(n669), .Z(n153) );
  OR2 C6303 ( .A(n153), .B(n726), .Z(n152) );
  OR2 C6302 ( .A(n152), .B(n781), .Z(n151) );
  OR2 C6301 ( .A(n151), .B(n888), .Z(n150) );
  AN2 C6300 ( .A(ENCODER_CONTROL_IN[6]), .B(n150), .Z(n1783) );
  OR2 C6298 ( .A(n412), .B(n470), .Z(n163) );
  OR2 C6297 ( .A(n163), .B(n593), .Z(n162) );
  OR2 C6296 ( .A(n162), .B(n534), .Z(n161) );
  OR2 C6295 ( .A(n161), .B(n654), .Z(n160) );
  OR2 C6294 ( .A(n160), .B(n713), .Z(n159) );
  OR2 C6293 ( .A(n159), .B(n764), .Z(n158) );
  OR2 C6292 ( .A(n158), .B(n873), .Z(n157) );
  AN2 C6291 ( .A(ENCODER_CONTROL_IN[5]), .B(n157), .Z(n1785) );
  OR2 C6289 ( .A(n405), .B(n463), .Z(n170) );
  OR2 C6288 ( .A(n170), .B(n586), .Z(n169) );
  OR2 C6287 ( .A(n169), .B(n526), .Z(n168) );
  OR2 C6286 ( .A(n168), .B(n646), .Z(n167) );
  OR2 C6285 ( .A(n167), .B(n706), .Z(n166) );
  OR2 C6284 ( .A(n166), .B(n758), .Z(n165) );
  OR2 C6283 ( .A(n165), .B(n862), .Z(n164) );
  AN2 C6282 ( .A(ENCODER_CONTROL_IN[4]), .B(n164), .Z(n1787) );
  OR2 C6280 ( .A(n398), .B(n455), .Z(n177) );
  OR2 C6279 ( .A(n177), .B(n579), .Z(n176) );
  OR2 C6278 ( .A(n176), .B(n518), .Z(n175) );
  OR2 C6277 ( .A(n175), .B(n638), .Z(n174) );
  OR2 C6276 ( .A(n174), .B(n699), .Z(n173) );
  OR2 C6275 ( .A(n173), .B(n752), .Z(n172) );
  OR2 C6274 ( .A(n172), .B(n823), .Z(n171) );
  AN2 C6273 ( .A(ENCODER_CONTROL_IN[3]), .B(n171), .Z(n1789) );
  OR2 C6271 ( .A(n391), .B(n447), .Z(n184) );
  OR2 C6270 ( .A(n184), .B(n572), .Z(n183) );
  OR2 C6269 ( .A(n183), .B(n510), .Z(n182) );
  OR2 C6268 ( .A(n182), .B(n630), .Z(n181) );
  OR2 C6267 ( .A(n181), .B(n692), .Z(n180) );
  OR2 C6266 ( .A(n180), .B(n746), .Z(n179) );
  OR2 C6265 ( .A(n179), .B(n808), .Z(n178) );
  AN2 C6264 ( .A(ENCODER_CONTROL_IN[2]), .B(n178), .Z(n1791) );
  OR2 C6262 ( .A(n384), .B(n432), .Z(n191) );
  OR2 C6261 ( .A(n191), .B(n557), .Z(n190) );
  OR2 C6260 ( .A(n190), .B(n494), .Z(n189) );
  OR2 C6259 ( .A(n189), .B(n615), .Z(n188) );
  OR2 C6258 ( .A(n188), .B(n677), .Z(n187) );
  OR2 C6257 ( .A(n187), .B(n733), .Z(n186) );
  OR2 C6256 ( .A(n186), .B(n787), .Z(n185) );
  AN2 C6255 ( .A(ENCODER_CONTROL_IN[1]), .B(n185), .Z(n1793) );
  OR2 C6253 ( .A(n377), .B(n418), .Z(n198) );
  OR2 C6252 ( .A(n198), .B(n542), .Z(n197) );
  OR2 C6251 ( .A(n197), .B(n478), .Z(n196) );
  OR2 C6250 ( .A(n196), .B(n600), .Z(n195) );
  OR2 C6249 ( .A(n195), .B(n662), .Z(n194) );
  OR2 C6248 ( .A(n194), .B(n720), .Z(n193) );
  OR2 C6247 ( .A(n193), .B(n770), .Z(n192) );
  AN2 C6246 ( .A(ENCODER_CONTROL_IN[0]), .B(n192), .Z(n1795) );
  AN2 C6244 ( .A(ENCODER_CONTROL_IN[4]), .B(n337), .Z(n1797) );
  AN2 C6242 ( .A(ENCODER_CONTROL_IN[0]), .B(n348), .Z(n1799) );
  AN2 C6240 ( .A(ENCODER_CONTROL_IN[4]), .B(n850), .Z(n1801) );
  OR2 C6238 ( .A(n330), .B(n850), .Z(n199) );
  AN2 C6237 ( .A(ENCODER_CONTROL_IN[4]), .B(n199), .Z(n1803) );
  AN2 C6235 ( .A(ENCODER_CONTROL_IN[0]), .B(n838), .Z(n1805) );
  OR2 C6233 ( .A(n341), .B(n838), .Z(n200) );
  AN2 C6232 ( .A(ENCODER_CONTROL_IN[0]), .B(n200), .Z(n1807) );
  AN2 C6230 ( .A(ENCODER_CONTROL_IN[7]), .B(n373), .Z(n1809) );
  AN2 C6228 ( .A(ENCODER_CONTROL_IN[6]), .B(n370), .Z(n1811) );
  AN2 C6226 ( .A(ENCODER_CONTROL_IN[5]), .B(n367), .Z(n1813) );
  AN2 C6224 ( .A(ENCODER_CONTROL_IN[4]), .B(n364), .Z(n1815) );
  AN2 C6222 ( .A(ENCODER_CONTROL_IN[3]), .B(n361), .Z(n1817) );
  AN2 C6220 ( .A(ENCODER_CONTROL_IN[2]), .B(n358), .Z(n1819) );
  AN2 C6218 ( .A(ENCODER_CONTROL_IN[1]), .B(n355), .Z(n1821) );
  AN2 C6216 ( .A(ENCODER_CONTROL_IN[0]), .B(n352), .Z(n1823) );
  AN2 C5895 ( .A(n1960), .B(ENCODER_CONTROL_IN[0]), .Z(n201) );
  AN2 C5894 ( .A(n1951), .B(ENCODER_CONTROL_IN[1]), .Z(n203) );
  AN2 C5893 ( .A(n1950), .B(ENCODER_CONTROL_IN[2]), .Z(n205) );
  AN2 C5892 ( .A(n1949), .B(ENCODER_CONTROL_IN[3]), .Z(n207) );
  AN2 C5891 ( .A(n1948), .B(ENCODER_CONTROL_IN[4]), .Z(n209) );
  AN2 C5890 ( .A(n1947), .B(ENCODER_CONTROL_IN[5]), .Z(n211) );
  AN2 C5889 ( .A(n1946), .B(ENCODER_CONTROL_IN[6]), .Z(n213) );
  AN2 C5888 ( .A(n1945), .B(ENCODER_CONTROL_IN[7]), .Z(n214) );
  OR2 C5887 ( .A(n214), .B(n213), .Z(n212) );
  OR2 C5886 ( .A(n212), .B(n211), .Z(n210) );
  OR2 C5885 ( .A(n210), .B(n209), .Z(n208) );
  OR2 C5884 ( .A(n208), .B(n207), .Z(n206) );
  OR2 C5883 ( .A(n206), .B(n205), .Z(n204) );
  OR2 C5882 ( .A(n204), .B(n203), .Z(n202) );
  OR2 C5881 ( .A(n202), .B(n201), .Z(n1944) );
  AN2 C5879 ( .A(n374), .B(n442), .Z(n221) );
  AN2 C5878 ( .A(n221), .B(n503), .Z(n220) );
  AN2 C5877 ( .A(n220), .B(n624), .Z(n219) );
  AN2 C5876 ( .A(n219), .B(n565), .Z(n218) );
  AN2 C5875 ( .A(n218), .B(n685), .Z(n217) );
  AN2 C5874 ( .A(n217), .B(n740), .Z(n216) );
  AN2 C5873 ( .A(n216), .B(n803), .Z(n215) );
  AN2 C5872 ( .A(n215), .B(n904), .Z(n1945) );
  AN2 C5870 ( .A(n371), .B(n427), .Z(n228) );
  AN2 C5869 ( .A(n228), .B(n487), .Z(n227) );
  AN2 C5868 ( .A(n227), .B(n609), .Z(n226) );
  AN2 C5867 ( .A(n226), .B(n550), .Z(n225) );
  AN2 C5866 ( .A(n225), .B(n670), .Z(n224) );
  AN2 C5865 ( .A(n224), .B(n727), .Z(n223) );
  AN2 C5864 ( .A(n223), .B(n782), .Z(n222) );
  AN2 C5863 ( .A(n222), .B(n889), .Z(n1946) );
  AN2 C5861 ( .A(n368), .B(n413), .Z(n235) );
  AN2 C5860 ( .A(n235), .B(n471), .Z(n234) );
  AN2 C5859 ( .A(n234), .B(n594), .Z(n233) );
  AN2 C5858 ( .A(n233), .B(n535), .Z(n232) );
  AN2 C5857 ( .A(n232), .B(n655), .Z(n231) );
  AN2 C5856 ( .A(n231), .B(n714), .Z(n230) );
  AN2 C5855 ( .A(n230), .B(n765), .Z(n229) );
  AN2 C5854 ( .A(n229), .B(n874), .Z(n1947) );
  AN2 C5852 ( .A(n365), .B(n851), .Z(n245) );
  AN2 C5851 ( .A(n245), .B(n338), .Z(n244) );
  AN2 C5850 ( .A(n244), .B(n331), .Z(n243) );
  AN2 C5849 ( .A(n243), .B(n406), .Z(n242) );
  AN2 C5848 ( .A(n242), .B(n464), .Z(n241) );
  AN2 C5847 ( .A(n241), .B(n587), .Z(n240) );
  AN2 C5846 ( .A(n240), .B(n527), .Z(n239) );
  AN2 C5845 ( .A(n239), .B(n647), .Z(n238) );
  AN2 C5844 ( .A(n238), .B(n707), .Z(n237) );
  AN2 C5843 ( .A(n237), .B(n759), .Z(n236) );
  AN2 C5842 ( .A(n236), .B(n863), .Z(n1948) );
  AN2 C5840 ( .A(n362), .B(n399), .Z(n252) );
  AN2 C5839 ( .A(n252), .B(n456), .Z(n251) );
  AN2 C5838 ( .A(n251), .B(n580), .Z(n250) );
  AN2 C5837 ( .A(n250), .B(n519), .Z(n249) );
  AN2 C5836 ( .A(n249), .B(n639), .Z(n248) );
  AN2 C5835 ( .A(n248), .B(n700), .Z(n247) );
  AN2 C5834 ( .A(n247), .B(n753), .Z(n246) );
  AN2 C5833 ( .A(n246), .B(n824), .Z(n1949) );
  AN2 C5831 ( .A(n359), .B(n392), .Z(n259) );
  AN2 C5830 ( .A(n259), .B(n448), .Z(n258) );
  AN2 C5829 ( .A(n258), .B(n573), .Z(n257) );
  AN2 C5828 ( .A(n257), .B(n511), .Z(n256) );
  AN2 C5827 ( .A(n256), .B(n631), .Z(n255) );
  AN2 C5826 ( .A(n255), .B(n693), .Z(n254) );
  AN2 C5825 ( .A(n254), .B(n747), .Z(n253) );
  AN2 C5824 ( .A(n253), .B(n809), .Z(n1950) );
  AN2 C5822 ( .A(n356), .B(n385), .Z(n266) );
  AN2 C5821 ( .A(n266), .B(n433), .Z(n265) );
  AN2 C5820 ( .A(n265), .B(n558), .Z(n264) );
  AN2 C5819 ( .A(n264), .B(n495), .Z(n263) );
  AN2 C5818 ( .A(n263), .B(n616), .Z(n262) );
  AN2 C5817 ( .A(n262), .B(n678), .Z(n261) );
  AN2 C5816 ( .A(n261), .B(n734), .Z(n260) );
  AN2 C5815 ( .A(n260), .B(n788), .Z(n1951) );
  AN2 C5813 ( .A(n353), .B(n839), .Z(n276) );
  AN2 C5812 ( .A(n276), .B(n349), .Z(n275) );
  AN2 C5811 ( .A(n275), .B(n342), .Z(n274) );
  AN2 C5810 ( .A(n274), .B(n378), .Z(n273) );
  AN2 C5809 ( .A(n273), .B(n419), .Z(n272) );
  AN2 C5808 ( .A(n272), .B(n543), .Z(n271) );
  AN2 C5807 ( .A(n271), .B(n479), .Z(n270) );
  AN2 C5806 ( .A(n270), .B(n601), .Z(n269) );
  AN2 C5805 ( .A(n269), .B(n663), .Z(n268) );
  AN2 C5804 ( .A(n268), .B(n721), .Z(n267) );
  AN2 C5803 ( .A(n267), .B(n771), .Z(n1960) );
  IV I_170 ( .A(ENCODER_CONTROL_IN[7]), .Z(n1961) );
  IV I_169 ( .A(ENCODER_CONTROL_IN[6]), .Z(n1962) );
  IV I_168 ( .A(ENCODER_CONTROL_IN[5]), .Z(n1963) );
  IV I_167 ( .A(ENCODER_CONTROL_IN[4]), .Z(n1964) );
  IV I_166 ( .A(ENCODER_CONTROL_IN[3]), .Z(n1965) );
  IV I_165 ( .A(ENCODER_CONTROL_IN[2]), .Z(n1966) );
  IV I_164 ( .A(ENCODER_CONTROL_IN[1]), .Z(n1967) );
  IV I_163 ( .A(ENCODER_CONTROL_IN[0]), .Z(n1968) );
  AN2 C5792 ( .A(n2491), .B(n959), .Z(ENCODER_DATA_OUT[1]) );
  OR2 C5646 ( .A(n1062), .B(n1237), .Z(n278) );
  OR2 C5458 ( .A(n1297), .B(n1363), .Z(n279) );
  OR2 C5455 ( .A(n1297), .B(n1296), .Z(n281) );
  OR2 C5421 ( .A(n297), .B(n284), .Z(n283) );
  OR2 C5379 ( .A(n297), .B(n287), .Z(n286) );
  OR2 C5335 ( .A(n297), .B(n290), .Z(n289) );
  OR2 C5334 ( .A(n1503), .B(n1487), .Z(n290) );
  OR2 C5294 ( .A(n1647), .B(n1599), .Z(n295) );
  OR2 C5293 ( .A(n297), .B(n1503), .Z(n296) );
  OR2 C5256 ( .A(U29_CONTROL1), .B(n1519), .Z(n301) );
  OR2 C5194 ( .A(n306), .B(n1439), .Z(n305) );
  OR2 C5145 ( .A(n310), .B(n309), .Z(n308) );
  OR2 C5144 ( .A(n1455), .B(n1439), .Z(n309) );
  OR2 C5138 ( .A(n314), .B(U19_CONTROL4), .Z(U10_DATA2_7) );
  OR2 C5131 ( .A(n316), .B(U19_CONTROL4), .Z(U10_DATA2_6) );
  OR2 C5124 ( .A(n319), .B(n318), .Z(U10_DATA2_5) );
  OR2 C5114 ( .A(n321), .B(n320), .Z(U10_DATA2_4) );
  OR2 C5107 ( .A(n323), .B(n322), .Z(U10_DATA2_3) );
  OR2 C5100 ( .A(n325), .B(n324), .Z(U10_DATA2_2) );
  OR2 C5093 ( .A(n327), .B(n326), .Z(U10_DATA2_1) );
  OR2 C5089 ( .A(n329), .B(n328), .Z(U10_DATA2_0) );
  IV I_160 ( .A(n331), .Z(n330) );
  OR2 C2879 ( .A(ENCODER_DATA_IN[32]), .B(n332), .Z(n331) );
  OR2 C2878 ( .A(ENCODER_DATA_IN[33]), .B(n333), .Z(n332) );
  OR2 C2877 ( .A(n858), .B(n334), .Z(n333) );
  OR2 C2876 ( .A(n859), .B(n335), .Z(n334) );
  OR2 C2875 ( .A(n860), .B(n336), .Z(n335) );
  OR2 C2874 ( .A(ENCODER_DATA_IN[37]), .B(n533), .Z(n336) );
  IV I_159 ( .A(n338), .Z(n337) );
  OR2 C2867 ( .A(n763), .B(n339), .Z(n338) );
  OR2 C2866 ( .A(n870), .B(n340), .Z(n339) );
  OR2 C2865 ( .A(ENCODER_DATA_IN[34]), .B(n866), .Z(n340) );
  IV I_158 ( .A(n342), .Z(n341) );
  OR2 C2840 ( .A(ENCODER_DATA_IN[0]), .B(n343), .Z(n342) );
  OR2 C2839 ( .A(ENCODER_DATA_IN[1]), .B(n344), .Z(n343) );
  OR2 C2838 ( .A(n846), .B(n345), .Z(n344) );
  OR2 C2837 ( .A(n847), .B(n346), .Z(n345) );
  OR2 C2836 ( .A(n848), .B(n347), .Z(n346) );
  OR2 C2835 ( .A(ENCODER_DATA_IN[5]), .B(n485), .Z(n347) );
  IV I_157 ( .A(n349), .Z(n348) );
  OR2 C2828 ( .A(n725), .B(n350), .Z(n349) );
  OR2 C2827 ( .A(n778), .B(n351), .Z(n350) );
  OR2 C2826 ( .A(ENCODER_DATA_IN[2]), .B(n774), .Z(n351) );
  IV I_156 ( .A(n353), .Z(n352) );
  OR2 C2813 ( .A(n725), .B(n354), .Z(n353) );
  OR2 C2812 ( .A(ENCODER_DATA_IN[1]), .B(n773), .Z(n354) );
  IV I_155 ( .A(n356), .Z(n355) );
  OR2 C2798 ( .A(n738), .B(n357), .Z(n356) );
  OR2 C2797 ( .A(ENCODER_DATA_IN[9]), .B(n790), .Z(n357) );
  IV I_154 ( .A(n359), .Z(n358) );
  OR2 C2783 ( .A(n751), .B(n360), .Z(n359) );
  OR2 C2782 ( .A(ENCODER_DATA_IN[17]), .B(n811), .Z(n360) );
  IV I_153 ( .A(n362), .Z(n361) );
  OR2 C2768 ( .A(n757), .B(n363), .Z(n362) );
  OR2 C2767 ( .A(ENCODER_DATA_IN[25]), .B(n826), .Z(n363) );
  IV I_152 ( .A(n365), .Z(n364) );
  OR2 C2753 ( .A(n763), .B(n366), .Z(n365) );
  OR2 C2752 ( .A(ENCODER_DATA_IN[33]), .B(n865), .Z(n366) );
  IV I_151 ( .A(n368), .Z(n367) );
  OR2 C2738 ( .A(n769), .B(n369), .Z(n368) );
  OR2 C2737 ( .A(ENCODER_DATA_IN[41]), .B(n876), .Z(n369) );
  IV I_150 ( .A(n371), .Z(n370) );
  OR2 C2723 ( .A(n786), .B(n372), .Z(n371) );
  OR2 C2722 ( .A(ENCODER_DATA_IN[49]), .B(n891), .Z(n372) );
  IV I_149 ( .A(n374), .Z(n373) );
  OR2 C2708 ( .A(n807), .B(n375), .Z(n374) );
  OR2 C2707 ( .A(ENCODER_DATA_IN[57]), .B(n906), .Z(n375) );
  IV I_148 ( .A(ENCODER_CONTROL_IN[0]), .Z(n376) );
  IV I_147 ( .A(n378), .Z(n377) );
  OR2 C2692 ( .A(n725), .B(n379), .Z(n378) );
  OR2 C2691 ( .A(n778), .B(n380), .Z(n379) );
  OR2 C2690 ( .A(n846), .B(n381), .Z(n380) );
  OR2 C2689 ( .A(ENCODER_DATA_IN[3]), .B(n382), .Z(n381) );
  OR2 C2688 ( .A(ENCODER_DATA_IN[4]), .B(n548), .Z(n382) );
  IV I_146 ( .A(ENCODER_CONTROL_IN[1]), .Z(n383) );
  IV I_145 ( .A(n385), .Z(n384) );
  OR2 C2680 ( .A(n738), .B(n386), .Z(n385) );
  OR2 C2679 ( .A(n795), .B(n387), .Z(n386) );
  OR2 C2678 ( .A(n796), .B(n388), .Z(n387) );
  OR2 C2677 ( .A(ENCODER_DATA_IN[11]), .B(n389), .Z(n388) );
  OR2 C2676 ( .A(ENCODER_DATA_IN[12]), .B(n563), .Z(n389) );
  IV I_144 ( .A(ENCODER_CONTROL_IN[2]), .Z(n390) );
  IV I_143 ( .A(n392), .Z(n391) );
  OR2 C2668 ( .A(n751), .B(n393), .Z(n392) );
  OR2 C2667 ( .A(n816), .B(n394), .Z(n393) );
  OR2 C2666 ( .A(n817), .B(n395), .Z(n394) );
  OR2 C2665 ( .A(ENCODER_DATA_IN[19]), .B(n396), .Z(n395) );
  OR2 C2664 ( .A(ENCODER_DATA_IN[20]), .B(n578), .Z(n396) );
  IV I_142 ( .A(ENCODER_CONTROL_IN[3]), .Z(n397) );
  IV I_141 ( .A(n399), .Z(n398) );
  OR2 C2656 ( .A(n757), .B(n400), .Z(n399) );
  OR2 C2655 ( .A(n831), .B(n401), .Z(n400) );
  OR2 C2654 ( .A(n832), .B(n402), .Z(n401) );
  OR2 C2653 ( .A(ENCODER_DATA_IN[27]), .B(n403), .Z(n402) );
  OR2 C2652 ( .A(ENCODER_DATA_IN[28]), .B(n585), .Z(n403) );
  IV I_140 ( .A(ENCODER_CONTROL_IN[4]), .Z(n404) );
  IV I_139 ( .A(n406), .Z(n405) );
  OR2 C2644 ( .A(n763), .B(n407), .Z(n406) );
  OR2 C2643 ( .A(n870), .B(n408), .Z(n407) );
  OR2 C2642 ( .A(n858), .B(n409), .Z(n408) );
  OR2 C2641 ( .A(ENCODER_DATA_IN[35]), .B(n410), .Z(n409) );
  OR2 C2640 ( .A(ENCODER_DATA_IN[36]), .B(n592), .Z(n410) );
  IV I_138 ( .A(ENCODER_CONTROL_IN[5]), .Z(n411) );
  IV I_137 ( .A(n413), .Z(n412) );
  OR2 C2632 ( .A(n769), .B(n414), .Z(n413) );
  OR2 C2631 ( .A(n881), .B(n415), .Z(n414) );
  OR2 C2630 ( .A(n882), .B(n416), .Z(n415) );
  OR2 C2629 ( .A(ENCODER_DATA_IN[43]), .B(n417), .Z(n416) );
  OR2 C2628 ( .A(ENCODER_DATA_IN[44]), .B(n599), .Z(n417) );
  IV I_136 ( .A(n419), .Z(n418) );
  OR2 C2621 ( .A(ENCODER_DATA_IN[0]), .B(n420), .Z(n419) );
  OR2 C2620 ( .A(ENCODER_DATA_IN[1]), .B(n421), .Z(n420) );
  OR2 C2619 ( .A(n846), .B(n422), .Z(n421) );
  OR2 C2618 ( .A(n847), .B(n423), .Z(n422) );
  OR2 C2617 ( .A(n848), .B(n424), .Z(n423) );
  OR2 C2616 ( .A(n779), .B(n845), .Z(n424) );
  IV I_135 ( .A(ENCODER_CONTROL_IN[6]), .Z(n425) );
  IV I_134 ( .A(n427), .Z(n426) );
  OR2 C2607 ( .A(n786), .B(n428), .Z(n427) );
  OR2 C2606 ( .A(n896), .B(n429), .Z(n428) );
  OR2 C2605 ( .A(n897), .B(n430), .Z(n429) );
  OR2 C2604 ( .A(ENCODER_DATA_IN[51]), .B(n431), .Z(n430) );
  OR2 C2603 ( .A(ENCODER_DATA_IN[52]), .B(n614), .Z(n431) );
  IV I_133 ( .A(n433), .Z(n432) );
  OR2 C2596 ( .A(ENCODER_DATA_IN[8]), .B(n434), .Z(n433) );
  OR2 C2595 ( .A(ENCODER_DATA_IN[9]), .B(n435), .Z(n434) );
  OR2 C2594 ( .A(n796), .B(n436), .Z(n435) );
  OR2 C2593 ( .A(n797), .B(n437), .Z(n436) );
  OR2 C2592 ( .A(n798), .B(n438), .Z(n437) );
  OR2 C2591 ( .A(n799), .B(n439), .Z(n438) );
  OR2 C2590 ( .A(n800), .B(ENCODER_DATA_IN[15]), .Z(n439) );
  IV I_132 ( .A(ENCODER_CONTROL_IN[7]), .Z(n440) );
  IV I_131 ( .A(n442), .Z(n441) );
  OR2 C2582 ( .A(n807), .B(n443), .Z(n442) );
  OR2 C2581 ( .A(n911), .B(n444), .Z(n443) );
  OR2 C2580 ( .A(n912), .B(n445), .Z(n444) );
  OR2 C2579 ( .A(ENCODER_DATA_IN[59]), .B(n446), .Z(n445) );
  OR2 C2578 ( .A(ENCODER_DATA_IN[60]), .B(n629), .Z(n446) );
  IV I_130 ( .A(n448), .Z(n447) );
  OR2 C2571 ( .A(ENCODER_DATA_IN[16]), .B(n449), .Z(n448) );
  OR2 C2570 ( .A(ENCODER_DATA_IN[17]), .B(n450), .Z(n449) );
  OR2 C2569 ( .A(n817), .B(n451), .Z(n450) );
  OR2 C2568 ( .A(n818), .B(n452), .Z(n451) );
  OR2 C2567 ( .A(n819), .B(n453), .Z(n452) );
  OR2 C2566 ( .A(n820), .B(n454), .Z(n453) );
  OR2 C2565 ( .A(n821), .B(ENCODER_DATA_IN[23]), .Z(n454) );
  IV I_129 ( .A(n456), .Z(n455) );
  OR2 C2558 ( .A(ENCODER_DATA_IN[24]), .B(n457), .Z(n456) );
  OR2 C2557 ( .A(ENCODER_DATA_IN[25]), .B(n458), .Z(n457) );
  OR2 C2556 ( .A(n832), .B(n459), .Z(n458) );
  OR2 C2555 ( .A(n833), .B(n460), .Z(n459) );
  OR2 C2554 ( .A(n834), .B(n461), .Z(n460) );
  OR2 C2553 ( .A(n835), .B(n462), .Z(n461) );
  OR2 C2552 ( .A(n836), .B(ENCODER_DATA_IN[31]), .Z(n462) );
  IV I_128 ( .A(n464), .Z(n463) );
  OR2 C2545 ( .A(ENCODER_DATA_IN[32]), .B(n465), .Z(n464) );
  OR2 C2544 ( .A(ENCODER_DATA_IN[33]), .B(n466), .Z(n465) );
  OR2 C2543 ( .A(n858), .B(n467), .Z(n466) );
  OR2 C2542 ( .A(n859), .B(n468), .Z(n467) );
  OR2 C2541 ( .A(n860), .B(n469), .Z(n468) );
  OR2 C2540 ( .A(n871), .B(n857), .Z(n469) );
  IV I_127 ( .A(n471), .Z(n470) );
  OR2 C2532 ( .A(ENCODER_DATA_IN[40]), .B(n472), .Z(n471) );
  OR2 C2531 ( .A(ENCODER_DATA_IN[41]), .B(n473), .Z(n472) );
  OR2 C2530 ( .A(n882), .B(n474), .Z(n473) );
  OR2 C2529 ( .A(n883), .B(n475), .Z(n474) );
  OR2 C2528 ( .A(n884), .B(n476), .Z(n475) );
  OR2 C2527 ( .A(n885), .B(n477), .Z(n476) );
  OR2 C2526 ( .A(n886), .B(ENCODER_DATA_IN[47]), .Z(n477) );
  IV I_126 ( .A(n479), .Z(n478) );
  OR2 C2519 ( .A(ENCODER_DATA_IN[0]), .B(n480), .Z(n479) );
  OR2 C2518 ( .A(ENCODER_DATA_IN[1]), .B(n481), .Z(n480) );
  OR2 C2517 ( .A(n846), .B(n482), .Z(n481) );
  OR2 C2516 ( .A(n847), .B(n483), .Z(n482) );
  OR2 C2515 ( .A(n848), .B(n484), .Z(n483) );
  OR2 C2514 ( .A(n779), .B(n485), .Z(n484) );
  OR2 C2513 ( .A(ENCODER_DATA_IN[6]), .B(n780), .Z(n485) );
  IV I_125 ( .A(n487), .Z(n486) );
  OR2 C2506 ( .A(ENCODER_DATA_IN[48]), .B(n488), .Z(n487) );
  OR2 C2505 ( .A(ENCODER_DATA_IN[49]), .B(n489), .Z(n488) );
  OR2 C2504 ( .A(n897), .B(n490), .Z(n489) );
  OR2 C2503 ( .A(n898), .B(n491), .Z(n490) );
  OR2 C2502 ( .A(n899), .B(n492), .Z(n491) );
  OR2 C2501 ( .A(n900), .B(n493), .Z(n492) );
  OR2 C2500 ( .A(n901), .B(ENCODER_DATA_IN[55]), .Z(n493) );
  IV I_124 ( .A(n495), .Z(n494) );
  OR2 C2493 ( .A(ENCODER_DATA_IN[8]), .B(n496), .Z(n495) );
  OR2 C2492 ( .A(ENCODER_DATA_IN[9]), .B(n497), .Z(n496) );
  OR2 C2491 ( .A(n796), .B(n498), .Z(n497) );
  OR2 C2490 ( .A(n797), .B(n499), .Z(n498) );
  OR2 C2489 ( .A(n798), .B(n500), .Z(n499) );
  OR2 C2488 ( .A(n799), .B(n501), .Z(n500) );
  OR2 C2487 ( .A(ENCODER_DATA_IN[14]), .B(n801), .Z(n501) );
  IV I_123 ( .A(n503), .Z(n502) );
  OR2 C2480 ( .A(ENCODER_DATA_IN[56]), .B(n504), .Z(n503) );
  OR2 C2479 ( .A(ENCODER_DATA_IN[57]), .B(n505), .Z(n504) );
  OR2 C2478 ( .A(n912), .B(n506), .Z(n505) );
  OR2 C2477 ( .A(n913), .B(n507), .Z(n506) );
  OR2 C2476 ( .A(n914), .B(n508), .Z(n507) );
  OR2 C2475 ( .A(n915), .B(n509), .Z(n508) );
  OR2 C2474 ( .A(n916), .B(ENCODER_DATA_IN[63]), .Z(n509) );
  IV I_122 ( .A(n511), .Z(n510) );
  OR2 C2467 ( .A(ENCODER_DATA_IN[16]), .B(n512), .Z(n511) );
  OR2 C2466 ( .A(ENCODER_DATA_IN[17]), .B(n513), .Z(n512) );
  OR2 C2465 ( .A(n817), .B(n514), .Z(n513) );
  OR2 C2464 ( .A(n818), .B(n515), .Z(n514) );
  OR2 C2463 ( .A(n819), .B(n516), .Z(n515) );
  OR2 C2462 ( .A(n820), .B(n517), .Z(n516) );
  OR2 C2461 ( .A(ENCODER_DATA_IN[22]), .B(n822), .Z(n517) );
  IV I_121 ( .A(n519), .Z(n518) );
  OR2 C2454 ( .A(ENCODER_DATA_IN[24]), .B(n520), .Z(n519) );
  OR2 C2453 ( .A(ENCODER_DATA_IN[25]), .B(n521), .Z(n520) );
  OR2 C2452 ( .A(n832), .B(n522), .Z(n521) );
  OR2 C2451 ( .A(n833), .B(n523), .Z(n522) );
  OR2 C2450 ( .A(n834), .B(n524), .Z(n523) );
  OR2 C2449 ( .A(n835), .B(n525), .Z(n524) );
  OR2 C2448 ( .A(ENCODER_DATA_IN[30]), .B(n837), .Z(n525) );
  IV I_120 ( .A(n527), .Z(n526) );
  OR2 C2441 ( .A(ENCODER_DATA_IN[32]), .B(n528), .Z(n527) );
  OR2 C2440 ( .A(ENCODER_DATA_IN[33]), .B(n529), .Z(n528) );
  OR2 C2439 ( .A(n858), .B(n530), .Z(n529) );
  OR2 C2438 ( .A(n859), .B(n531), .Z(n530) );
  OR2 C2437 ( .A(n860), .B(n532), .Z(n531) );
  OR2 C2436 ( .A(n871), .B(n533), .Z(n532) );
  OR2 C2435 ( .A(ENCODER_DATA_IN[38]), .B(n872), .Z(n533) );
  IV I_119 ( .A(n535), .Z(n534) );
  OR2 C2428 ( .A(ENCODER_DATA_IN[40]), .B(n536), .Z(n535) );
  OR2 C2427 ( .A(ENCODER_DATA_IN[41]), .B(n537), .Z(n536) );
  OR2 C2426 ( .A(n882), .B(n538), .Z(n537) );
  OR2 C2425 ( .A(n883), .B(n539), .Z(n538) );
  OR2 C2424 ( .A(n884), .B(n540), .Z(n539) );
  OR2 C2423 ( .A(n885), .B(n541), .Z(n540) );
  OR2 C2422 ( .A(ENCODER_DATA_IN[46]), .B(n887), .Z(n541) );
  IV I_118 ( .A(n543), .Z(n542) );
  OR2 C2415 ( .A(ENCODER_DATA_IN[0]), .B(n544), .Z(n543) );
  OR2 C2414 ( .A(ENCODER_DATA_IN[1]), .B(n545), .Z(n544) );
  OR2 C2413 ( .A(n846), .B(n546), .Z(n545) );
  OR2 C2412 ( .A(n847), .B(n547), .Z(n546) );
  OR2 C2411 ( .A(n848), .B(n548), .Z(n547) );
  OR2 C2410 ( .A(ENCODER_DATA_IN[5]), .B(n607), .Z(n548) );
  IV I_117 ( .A(n550), .Z(n549) );
  OR2 C2404 ( .A(ENCODER_DATA_IN[48]), .B(n551), .Z(n550) );
  OR2 C2403 ( .A(ENCODER_DATA_IN[49]), .B(n552), .Z(n551) );
  OR2 C2402 ( .A(n897), .B(n553), .Z(n552) );
  OR2 C2401 ( .A(n898), .B(n554), .Z(n553) );
  OR2 C2400 ( .A(n899), .B(n555), .Z(n554) );
  OR2 C2399 ( .A(n900), .B(n556), .Z(n555) );
  OR2 C2398 ( .A(ENCODER_DATA_IN[54]), .B(n902), .Z(n556) );
  IV I_116 ( .A(n558), .Z(n557) );
  OR2 C2391 ( .A(ENCODER_DATA_IN[8]), .B(n559), .Z(n558) );
  OR2 C2390 ( .A(ENCODER_DATA_IN[9]), .B(n560), .Z(n559) );
  OR2 C2389 ( .A(n796), .B(n561), .Z(n560) );
  OR2 C2388 ( .A(n797), .B(n562), .Z(n561) );
  OR2 C2387 ( .A(n798), .B(n563), .Z(n562) );
  OR2 C2386 ( .A(ENCODER_DATA_IN[13]), .B(n622), .Z(n563) );
  IV I_115 ( .A(n565), .Z(n564) );
  OR2 C2380 ( .A(ENCODER_DATA_IN[56]), .B(n566), .Z(n565) );
  OR2 C2379 ( .A(ENCODER_DATA_IN[57]), .B(n567), .Z(n566) );
  OR2 C2378 ( .A(n912), .B(n568), .Z(n567) );
  OR2 C2377 ( .A(n913), .B(n569), .Z(n568) );
  OR2 C2376 ( .A(n914), .B(n570), .Z(n569) );
  OR2 C2375 ( .A(n915), .B(n571), .Z(n570) );
  OR2 C2374 ( .A(ENCODER_DATA_IN[62]), .B(n917), .Z(n571) );
  IV I_114 ( .A(n573), .Z(n572) );
  OR2 C2367 ( .A(ENCODER_DATA_IN[16]), .B(n574), .Z(n573) );
  OR2 C2366 ( .A(ENCODER_DATA_IN[17]), .B(n575), .Z(n574) );
  OR2 C2365 ( .A(n817), .B(n576), .Z(n575) );
  OR2 C2364 ( .A(n818), .B(n577), .Z(n576) );
  OR2 C2363 ( .A(n819), .B(n578), .Z(n577) );
  OR2 C2362 ( .A(ENCODER_DATA_IN[21]), .B(n637), .Z(n578) );
  IV I_113 ( .A(n580), .Z(n579) );
  OR2 C2356 ( .A(ENCODER_DATA_IN[24]), .B(n581), .Z(n580) );
  OR2 C2355 ( .A(ENCODER_DATA_IN[25]), .B(n582), .Z(n581) );
  OR2 C2354 ( .A(n832), .B(n583), .Z(n582) );
  OR2 C2353 ( .A(n833), .B(n584), .Z(n583) );
  OR2 C2352 ( .A(n834), .B(n585), .Z(n584) );
  OR2 C2351 ( .A(ENCODER_DATA_IN[29]), .B(n645), .Z(n585) );
  IV I_112 ( .A(n587), .Z(n586) );
  OR2 C2345 ( .A(ENCODER_DATA_IN[32]), .B(n588), .Z(n587) );
  OR2 C2344 ( .A(ENCODER_DATA_IN[33]), .B(n589), .Z(n588) );
  OR2 C2343 ( .A(n858), .B(n590), .Z(n589) );
  OR2 C2342 ( .A(n859), .B(n591), .Z(n590) );
  OR2 C2341 ( .A(n860), .B(n592), .Z(n591) );
  OR2 C2340 ( .A(ENCODER_DATA_IN[37]), .B(n653), .Z(n592) );
  IV I_111 ( .A(n594), .Z(n593) );
  OR2 C2334 ( .A(ENCODER_DATA_IN[40]), .B(n595), .Z(n594) );
  OR2 C2333 ( .A(ENCODER_DATA_IN[41]), .B(n596), .Z(n595) );
  OR2 C2332 ( .A(n882), .B(n597), .Z(n596) );
  OR2 C2331 ( .A(n883), .B(n598), .Z(n597) );
  OR2 C2330 ( .A(n884), .B(n599), .Z(n598) );
  OR2 C2329 ( .A(ENCODER_DATA_IN[45]), .B(n661), .Z(n599) );
  IV I_110 ( .A(n601), .Z(n600) );
  OR2 C2323 ( .A(ENCODER_DATA_IN[0]), .B(n602), .Z(n601) );
  OR2 C2322 ( .A(ENCODER_DATA_IN[1]), .B(n603), .Z(n602) );
  OR2 C2321 ( .A(n846), .B(n604), .Z(n603) );
  OR2 C2320 ( .A(n847), .B(n605), .Z(n604) );
  OR2 C2319 ( .A(n848), .B(n606), .Z(n605) );
  OR2 C2318 ( .A(n779), .B(n607), .Z(n606) );
  OR2 C2317 ( .A(ENCODER_DATA_IN[6]), .B(ENCODER_DATA_IN[7]), .Z(n607) );
  IV I_109 ( .A(n609), .Z(n608) );
  OR2 C2311 ( .A(ENCODER_DATA_IN[48]), .B(n610), .Z(n609) );
  OR2 C2310 ( .A(ENCODER_DATA_IN[49]), .B(n611), .Z(n610) );
  OR2 C2309 ( .A(n897), .B(n612), .Z(n611) );
  OR2 C2308 ( .A(n898), .B(n613), .Z(n612) );
  OR2 C2307 ( .A(n899), .B(n614), .Z(n613) );
  OR2 C2306 ( .A(ENCODER_DATA_IN[53]), .B(n676), .Z(n614) );
  IV I_108 ( .A(n616), .Z(n615) );
  OR2 C2300 ( .A(ENCODER_DATA_IN[8]), .B(n617), .Z(n616) );
  OR2 C2299 ( .A(ENCODER_DATA_IN[9]), .B(n618), .Z(n617) );
  OR2 C2298 ( .A(n796), .B(n619), .Z(n618) );
  OR2 C2297 ( .A(n797), .B(n620), .Z(n619) );
  OR2 C2296 ( .A(n798), .B(n621), .Z(n620) );
  OR2 C2295 ( .A(n799), .B(n622), .Z(n621) );
  OR2 C2294 ( .A(ENCODER_DATA_IN[14]), .B(ENCODER_DATA_IN[15]), .Z(n622) );
  IV I_107 ( .A(n624), .Z(n623) );
  OR2 C2288 ( .A(ENCODER_DATA_IN[56]), .B(n625), .Z(n624) );
  OR2 C2287 ( .A(ENCODER_DATA_IN[57]), .B(n626), .Z(n625) );
  OR2 C2286 ( .A(n912), .B(n627), .Z(n626) );
  OR2 C2285 ( .A(n913), .B(n628), .Z(n627) );
  OR2 C2284 ( .A(n914), .B(n629), .Z(n628) );
  OR2 C2283 ( .A(ENCODER_DATA_IN[61]), .B(n691), .Z(n629) );
  IV I_106 ( .A(n631), .Z(n630) );
  OR2 C2277 ( .A(ENCODER_DATA_IN[16]), .B(n632), .Z(n631) );
  OR2 C2276 ( .A(ENCODER_DATA_IN[17]), .B(n633), .Z(n632) );
  OR2 C2275 ( .A(n817), .B(n634), .Z(n633) );
  OR2 C2274 ( .A(n818), .B(n635), .Z(n634) );
  OR2 C2273 ( .A(n819), .B(n636), .Z(n635) );
  OR2 C2272 ( .A(n820), .B(n637), .Z(n636) );
  OR2 C2271 ( .A(ENCODER_DATA_IN[22]), .B(ENCODER_DATA_IN[23]), .Z(n637) );
  IV I_105 ( .A(n639), .Z(n638) );
  OR2 C2265 ( .A(ENCODER_DATA_IN[24]), .B(n640), .Z(n639) );
  OR2 C2264 ( .A(ENCODER_DATA_IN[25]), .B(n641), .Z(n640) );
  OR2 C2263 ( .A(n832), .B(n642), .Z(n641) );
  OR2 C2262 ( .A(n833), .B(n643), .Z(n642) );
  OR2 C2261 ( .A(n834), .B(n644), .Z(n643) );
  OR2 C2260 ( .A(n835), .B(n645), .Z(n644) );
  OR2 C2259 ( .A(ENCODER_DATA_IN[30]), .B(ENCODER_DATA_IN[31]), .Z(n645) );
  IV I_104 ( .A(n647), .Z(n646) );
  OR2 C2253 ( .A(ENCODER_DATA_IN[32]), .B(n648), .Z(n647) );
  OR2 C2252 ( .A(ENCODER_DATA_IN[33]), .B(n649), .Z(n648) );
  OR2 C2251 ( .A(n858), .B(n650), .Z(n649) );
  OR2 C2250 ( .A(n859), .B(n651), .Z(n650) );
  OR2 C2249 ( .A(n860), .B(n652), .Z(n651) );
  OR2 C2248 ( .A(n871), .B(n653), .Z(n652) );
  OR2 C2247 ( .A(ENCODER_DATA_IN[38]), .B(ENCODER_DATA_IN[39]), .Z(n653) );
  IV I_103 ( .A(n655), .Z(n654) );
  OR2 C2233 ( .A(ENCODER_DATA_IN[40]), .B(n656), .Z(n655) );
  OR2 C2232 ( .A(ENCODER_DATA_IN[41]), .B(n657), .Z(n656) );
  OR2 C2231 ( .A(n882), .B(n658), .Z(n657) );
  OR2 C2230 ( .A(n883), .B(n659), .Z(n658) );
  OR2 C2229 ( .A(n884), .B(n660), .Z(n659) );
  OR2 C2228 ( .A(n885), .B(n661), .Z(n660) );
  OR2 C2227 ( .A(ENCODER_DATA_IN[46]), .B(ENCODER_DATA_IN[47]), .Z(n661) );
  IV I_102 ( .A(n663), .Z(n662) );
  OR2 C2221 ( .A(ENCODER_DATA_IN[0]), .B(n664), .Z(n663) );
  OR2 C2220 ( .A(ENCODER_DATA_IN[1]), .B(n665), .Z(n664) );
  OR2 C2219 ( .A(n846), .B(n666), .Z(n665) );
  OR2 C2218 ( .A(n847), .B(n667), .Z(n666) );
  OR2 C2217 ( .A(n848), .B(n668), .Z(n667) );
  OR2 C2216 ( .A(ENCODER_DATA_IN[5]), .B(n777), .Z(n668) );
  IV I_101 ( .A(n670), .Z(n669) );
  OR2 C2208 ( .A(ENCODER_DATA_IN[48]), .B(n671), .Z(n670) );
  OR2 C2207 ( .A(ENCODER_DATA_IN[49]), .B(n672), .Z(n671) );
  OR2 C2206 ( .A(n897), .B(n673), .Z(n672) );
  OR2 C2205 ( .A(n898), .B(n674), .Z(n673) );
  OR2 C2204 ( .A(n899), .B(n675), .Z(n674) );
  OR2 C2203 ( .A(n900), .B(n676), .Z(n675) );
  OR2 C2202 ( .A(ENCODER_DATA_IN[54]), .B(ENCODER_DATA_IN[55]), .Z(n676) );
  IV I_100 ( .A(n678), .Z(n677) );
  OR2 C2196 ( .A(ENCODER_DATA_IN[8]), .B(n679), .Z(n678) );
  OR2 C2195 ( .A(ENCODER_DATA_IN[9]), .B(n680), .Z(n679) );
  OR2 C2194 ( .A(n796), .B(n681), .Z(n680) );
  OR2 C2193 ( .A(n797), .B(n682), .Z(n681) );
  OR2 C2192 ( .A(n798), .B(n683), .Z(n682) );
  OR2 C2191 ( .A(ENCODER_DATA_IN[13]), .B(n794), .Z(n683) );
  IV I_99 ( .A(n685), .Z(n684) );
  OR2 C2183 ( .A(ENCODER_DATA_IN[56]), .B(n686), .Z(n685) );
  OR2 C2182 ( .A(ENCODER_DATA_IN[57]), .B(n687), .Z(n686) );
  OR2 C2181 ( .A(n912), .B(n688), .Z(n687) );
  OR2 C2180 ( .A(n913), .B(n689), .Z(n688) );
  OR2 C2179 ( .A(n914), .B(n690), .Z(n689) );
  OR2 C2178 ( .A(n915), .B(n691), .Z(n690) );
  OR2 C2177 ( .A(ENCODER_DATA_IN[62]), .B(ENCODER_DATA_IN[63]), .Z(n691) );
  IV I_98 ( .A(n693), .Z(n692) );
  OR2 C2171 ( .A(ENCODER_DATA_IN[16]), .B(n694), .Z(n693) );
  OR2 C2170 ( .A(ENCODER_DATA_IN[17]), .B(n695), .Z(n694) );
  OR2 C2169 ( .A(n817), .B(n696), .Z(n695) );
  OR2 C2168 ( .A(n818), .B(n697), .Z(n696) );
  OR2 C2167 ( .A(n819), .B(n698), .Z(n697) );
  OR2 C2166 ( .A(ENCODER_DATA_IN[21]), .B(n815), .Z(n698) );
  IV I_97 ( .A(n700), .Z(n699) );
  OR2 C2158 ( .A(ENCODER_DATA_IN[24]), .B(n701), .Z(n700) );
  OR2 C2157 ( .A(ENCODER_DATA_IN[25]), .B(n702), .Z(n701) );
  OR2 C2156 ( .A(n832), .B(n703), .Z(n702) );
  OR2 C2155 ( .A(n833), .B(n704), .Z(n703) );
  OR2 C2154 ( .A(n834), .B(n705), .Z(n704) );
  OR2 C2153 ( .A(ENCODER_DATA_IN[29]), .B(n830), .Z(n705) );
  IV I_96 ( .A(n707), .Z(n706) );
  OR2 C2145 ( .A(ENCODER_DATA_IN[32]), .B(n708), .Z(n707) );
  OR2 C2144 ( .A(ENCODER_DATA_IN[33]), .B(n709), .Z(n708) );
  OR2 C2143 ( .A(n858), .B(n710), .Z(n709) );
  OR2 C2142 ( .A(n859), .B(n711), .Z(n710) );
  OR2 C2141 ( .A(n860), .B(n712), .Z(n711) );
  OR2 C2140 ( .A(ENCODER_DATA_IN[37]), .B(n869), .Z(n712) );
  IV I_95 ( .A(n714), .Z(n713) );
  OR2 C2132 ( .A(ENCODER_DATA_IN[40]), .B(n715), .Z(n714) );
  OR2 C2131 ( .A(ENCODER_DATA_IN[41]), .B(n716), .Z(n715) );
  OR2 C2130 ( .A(n882), .B(n717), .Z(n716) );
  OR2 C2129 ( .A(n883), .B(n718), .Z(n717) );
  OR2 C2128 ( .A(n884), .B(n719), .Z(n718) );
  OR2 C2127 ( .A(ENCODER_DATA_IN[45]), .B(n880), .Z(n719) );
  IV I_94 ( .A(n721), .Z(n720) );
  OR2 C2119 ( .A(n725), .B(n722), .Z(n721) );
  OR2 C2118 ( .A(n778), .B(n723), .Z(n722) );
  OR2 C2117 ( .A(n846), .B(n724), .Z(n723) );
  OR2 C2116 ( .A(ENCODER_DATA_IN[3]), .B(n775), .Z(n724) );
  IV I_93 ( .A(ENCODER_DATA_IN[0]), .Z(n725) );
  IV I_92 ( .A(n727), .Z(n726) );
  OR2 C2104 ( .A(ENCODER_DATA_IN[48]), .B(n728), .Z(n727) );
  OR2 C2103 ( .A(ENCODER_DATA_IN[49]), .B(n729), .Z(n728) );
  OR2 C2102 ( .A(n897), .B(n730), .Z(n729) );
  OR2 C2101 ( .A(n898), .B(n731), .Z(n730) );
  OR2 C2100 ( .A(n899), .B(n732), .Z(n731) );
  OR2 C2099 ( .A(ENCODER_DATA_IN[53]), .B(n895), .Z(n732) );
  IV I_91 ( .A(n734), .Z(n733) );
  OR2 C2091 ( .A(n738), .B(n735), .Z(n734) );
  OR2 C2090 ( .A(n795), .B(n736), .Z(n735) );
  OR2 C2089 ( .A(n796), .B(n737), .Z(n736) );
  OR2 C2088 ( .A(ENCODER_DATA_IN[11]), .B(n792), .Z(n737) );
  IV I_90 ( .A(ENCODER_DATA_IN[8]), .Z(n738) );
  IV I_89 ( .A(n740), .Z(n739) );
  OR2 C2076 ( .A(ENCODER_DATA_IN[56]), .B(n741), .Z(n740) );
  OR2 C2075 ( .A(ENCODER_DATA_IN[57]), .B(n742), .Z(n741) );
  OR2 C2074 ( .A(n912), .B(n743), .Z(n742) );
  OR2 C2073 ( .A(n913), .B(n744), .Z(n743) );
  OR2 C2072 ( .A(n914), .B(n745), .Z(n744) );
  OR2 C2071 ( .A(ENCODER_DATA_IN[61]), .B(n910), .Z(n745) );
  IV I_88 ( .A(n747), .Z(n746) );
  OR2 C2063 ( .A(n751), .B(n748), .Z(n747) );
  OR2 C2062 ( .A(n816), .B(n749), .Z(n748) );
  OR2 C2061 ( .A(n817), .B(n750), .Z(n749) );
  OR2 C2060 ( .A(ENCODER_DATA_IN[19]), .B(n813), .Z(n750) );
  IV I_87 ( .A(ENCODER_DATA_IN[16]), .Z(n751) );
  IV I_86 ( .A(n753), .Z(n752) );
  OR2 C2048 ( .A(n757), .B(n754), .Z(n753) );
  OR2 C2047 ( .A(n831), .B(n755), .Z(n754) );
  OR2 C2046 ( .A(n832), .B(n756), .Z(n755) );
  OR2 C2045 ( .A(ENCODER_DATA_IN[27]), .B(n828), .Z(n756) );
  IV I_85 ( .A(ENCODER_DATA_IN[24]), .Z(n757) );
  IV I_84 ( .A(n759), .Z(n758) );
  OR2 C2033 ( .A(n763), .B(n760), .Z(n759) );
  OR2 C2032 ( .A(n870), .B(n761), .Z(n760) );
  OR2 C2031 ( .A(n858), .B(n762), .Z(n761) );
  OR2 C2030 ( .A(ENCODER_DATA_IN[35]), .B(n867), .Z(n762) );
  IV I_83 ( .A(ENCODER_DATA_IN[32]), .Z(n763) );
  IV I_82 ( .A(n765), .Z(n764) );
  OR2 C2018 ( .A(n769), .B(n766), .Z(n765) );
  OR2 C2017 ( .A(n881), .B(n767), .Z(n766) );
  OR2 C2016 ( .A(n882), .B(n768), .Z(n767) );
  OR2 C2015 ( .A(ENCODER_DATA_IN[43]), .B(n878), .Z(n768) );
  IV I_81 ( .A(ENCODER_DATA_IN[40]), .Z(n769) );
  IV I_80 ( .A(n771), .Z(n770) );
  OR2 C2003 ( .A(ENCODER_DATA_IN[0]), .B(n772), .Z(n771) );
  OR2 C2002 ( .A(n778), .B(n773), .Z(n772) );
  OR2 C2001 ( .A(n846), .B(n774), .Z(n773) );
  OR2 C2000 ( .A(n847), .B(n775), .Z(n774) );
  OR2 C1999 ( .A(n848), .B(n776), .Z(n775) );
  OR2 C1998 ( .A(n779), .B(n777), .Z(n776) );
  OR2 C1997 ( .A(n849), .B(n780), .Z(n777) );
  IV I_79 ( .A(ENCODER_DATA_IN[1]), .Z(n778) );
  IV I_78 ( .A(ENCODER_DATA_IN[5]), .Z(n779) );
  IV I_77 ( .A(ENCODER_DATA_IN[7]), .Z(n780) );
  IV I_76 ( .A(n782), .Z(n781) );
  OR2 C1988 ( .A(n786), .B(n783), .Z(n782) );
  OR2 C1987 ( .A(n896), .B(n784), .Z(n783) );
  OR2 C1986 ( .A(n897), .B(n785), .Z(n784) );
  OR2 C1985 ( .A(ENCODER_DATA_IN[51]), .B(n893), .Z(n785) );
  IV I_75 ( .A(ENCODER_DATA_IN[48]), .Z(n786) );
  IV I_74 ( .A(n788), .Z(n787) );
  OR2 C1973 ( .A(ENCODER_DATA_IN[8]), .B(n789), .Z(n788) );
  OR2 C1972 ( .A(n795), .B(n790), .Z(n789) );
  OR2 C1971 ( .A(n796), .B(n791), .Z(n790) );
  OR2 C1970 ( .A(n797), .B(n792), .Z(n791) );
  OR2 C1969 ( .A(n798), .B(n793), .Z(n792) );
  OR2 C1968 ( .A(n799), .B(n794), .Z(n793) );
  OR2 C1967 ( .A(n800), .B(n801), .Z(n794) );
  IV I_73 ( .A(ENCODER_DATA_IN[9]), .Z(n795) );
  IV I_72 ( .A(ENCODER_DATA_IN[10]), .Z(n796) );
  IV I_71 ( .A(ENCODER_DATA_IN[11]), .Z(n797) );
  IV I_70 ( .A(ENCODER_DATA_IN[12]), .Z(n798) );
  IV I_69 ( .A(ENCODER_DATA_IN[13]), .Z(n799) );
  IV I_68 ( .A(ENCODER_DATA_IN[14]), .Z(n800) );
  IV I_67 ( .A(ENCODER_DATA_IN[15]), .Z(n801) );
  IV I_66 ( .A(n803), .Z(n802) );
  OR2 C1958 ( .A(n807), .B(n804), .Z(n803) );
  OR2 C1957 ( .A(n911), .B(n805), .Z(n804) );
  OR2 C1956 ( .A(n912), .B(n806), .Z(n805) );
  OR2 C1955 ( .A(ENCODER_DATA_IN[59]), .B(n908), .Z(n806) );
  IV I_65 ( .A(ENCODER_DATA_IN[56]), .Z(n807) );
  IV I_64 ( .A(n809), .Z(n808) );
  OR2 C1943 ( .A(ENCODER_DATA_IN[16]), .B(n810), .Z(n809) );
  OR2 C1942 ( .A(n816), .B(n811), .Z(n810) );
  OR2 C1941 ( .A(n817), .B(n812), .Z(n811) );
  OR2 C1940 ( .A(n818), .B(n813), .Z(n812) );
  OR2 C1939 ( .A(n819), .B(n814), .Z(n813) );
  OR2 C1938 ( .A(n820), .B(n815), .Z(n814) );
  OR2 C1937 ( .A(n821), .B(n822), .Z(n815) );
  IV I_63 ( .A(ENCODER_DATA_IN[17]), .Z(n816) );
  IV I_62 ( .A(ENCODER_DATA_IN[18]), .Z(n817) );
  IV I_61 ( .A(ENCODER_DATA_IN[19]), .Z(n818) );
  IV I_60 ( .A(ENCODER_DATA_IN[20]), .Z(n819) );
  IV I_59 ( .A(ENCODER_DATA_IN[21]), .Z(n820) );
  IV I_58 ( .A(ENCODER_DATA_IN[22]), .Z(n821) );
  IV I_57 ( .A(ENCODER_DATA_IN[23]), .Z(n822) );
  IV I_56 ( .A(n824), .Z(n823) );
  OR2 C1928 ( .A(ENCODER_DATA_IN[24]), .B(n825), .Z(n824) );
  OR2 C1927 ( .A(n831), .B(n826), .Z(n825) );
  OR2 C1926 ( .A(n832), .B(n827), .Z(n826) );
  OR2 C1925 ( .A(n833), .B(n828), .Z(n827) );
  OR2 C1924 ( .A(n834), .B(n829), .Z(n828) );
  OR2 C1923 ( .A(n835), .B(n830), .Z(n829) );
  OR2 C1922 ( .A(n836), .B(n837), .Z(n830) );
  IV I_55 ( .A(ENCODER_DATA_IN[25]), .Z(n831) );
  IV I_54 ( .A(ENCODER_DATA_IN[26]), .Z(n832) );
  IV I_53 ( .A(ENCODER_DATA_IN[27]), .Z(n833) );
  IV I_52 ( .A(ENCODER_DATA_IN[28]), .Z(n834) );
  IV I_51 ( .A(ENCODER_DATA_IN[29]), .Z(n835) );
  IV I_50 ( .A(ENCODER_DATA_IN[30]), .Z(n836) );
  IV I_49 ( .A(ENCODER_DATA_IN[31]), .Z(n837) );
  IV I_48 ( .A(n839), .Z(n838) );
  OR2 C1913 ( .A(ENCODER_DATA_IN[0]), .B(n840), .Z(n839) );
  OR2 C1912 ( .A(ENCODER_DATA_IN[1]), .B(n841), .Z(n840) );
  OR2 C1911 ( .A(n846), .B(n842), .Z(n841) );
  OR2 C1910 ( .A(n847), .B(n843), .Z(n842) );
  OR2 C1909 ( .A(n848), .B(n844), .Z(n843) );
  OR2 C1908 ( .A(ENCODER_DATA_IN[5]), .B(n845), .Z(n844) );
  OR2 C1907 ( .A(n849), .B(ENCODER_DATA_IN[7]), .Z(n845) );
  IV I_47 ( .A(ENCODER_DATA_IN[2]), .Z(n846) );
  IV I_46 ( .A(ENCODER_DATA_IN[3]), .Z(n847) );
  IV I_45 ( .A(ENCODER_DATA_IN[4]), .Z(n848) );
  IV I_44 ( .A(ENCODER_DATA_IN[6]), .Z(n849) );
  IV I_43 ( .A(n851), .Z(n850) );
  OR2 C1901 ( .A(ENCODER_DATA_IN[32]), .B(n852), .Z(n851) );
  OR2 C1900 ( .A(ENCODER_DATA_IN[33]), .B(n853), .Z(n852) );
  OR2 C1899 ( .A(n858), .B(n854), .Z(n853) );
  OR2 C1898 ( .A(n859), .B(n855), .Z(n854) );
  OR2 C1897 ( .A(n860), .B(n856), .Z(n855) );
  OR2 C1896 ( .A(ENCODER_DATA_IN[37]), .B(n857), .Z(n856) );
  OR2 C1895 ( .A(n861), .B(ENCODER_DATA_IN[39]), .Z(n857) );
  IV I_42 ( .A(ENCODER_DATA_IN[34]), .Z(n858) );
  IV I_41 ( .A(ENCODER_DATA_IN[35]), .Z(n859) );
  IV I_40 ( .A(ENCODER_DATA_IN[36]), .Z(n860) );
  IV I_39 ( .A(ENCODER_DATA_IN[38]), .Z(n861) );
  IV I_38 ( .A(n863), .Z(n862) );
  OR2 C1889 ( .A(ENCODER_DATA_IN[32]), .B(n864), .Z(n863) );
  OR2 C1888 ( .A(n870), .B(n865), .Z(n864) );
  OR2 C1887 ( .A(n858), .B(n866), .Z(n865) );
  OR2 C1886 ( .A(n859), .B(n867), .Z(n866) );
  OR2 C1885 ( .A(n860), .B(n868), .Z(n867) );
  OR2 C1884 ( .A(n871), .B(n869), .Z(n868) );
  OR2 C1883 ( .A(n861), .B(n872), .Z(n869) );
  IV I_37 ( .A(ENCODER_DATA_IN[33]), .Z(n870) );
  IV I_36 ( .A(ENCODER_DATA_IN[37]), .Z(n871) );
  IV I_35 ( .A(ENCODER_DATA_IN[39]), .Z(n872) );
  IV I_34 ( .A(n874), .Z(n873) );
  OR2 C1874 ( .A(ENCODER_DATA_IN[40]), .B(n875), .Z(n874) );
  OR2 C1873 ( .A(n881), .B(n876), .Z(n875) );
  OR2 C1872 ( .A(n882), .B(n877), .Z(n876) );
  OR2 C1871 ( .A(n883), .B(n878), .Z(n877) );
  OR2 C1870 ( .A(n884), .B(n879), .Z(n878) );
  OR2 C1869 ( .A(n885), .B(n880), .Z(n879) );
  OR2 C1868 ( .A(n886), .B(n887), .Z(n880) );
  IV I_33 ( .A(ENCODER_DATA_IN[41]), .Z(n881) );
  IV I_32 ( .A(ENCODER_DATA_IN[42]), .Z(n882) );
  IV I_31 ( .A(ENCODER_DATA_IN[43]), .Z(n883) );
  IV I_30 ( .A(ENCODER_DATA_IN[44]), .Z(n884) );
  IV I_29 ( .A(ENCODER_DATA_IN[45]), .Z(n885) );
  IV I_28 ( .A(ENCODER_DATA_IN[46]), .Z(n886) );
  IV I_27 ( .A(ENCODER_DATA_IN[47]), .Z(n887) );
  IV I_26 ( .A(n889), .Z(n888) );
  OR2 C1859 ( .A(ENCODER_DATA_IN[48]), .B(n890), .Z(n889) );
  OR2 C1858 ( .A(n896), .B(n891), .Z(n890) );
  OR2 C1857 ( .A(n897), .B(n892), .Z(n891) );
  OR2 C1856 ( .A(n898), .B(n893), .Z(n892) );
  OR2 C1855 ( .A(n899), .B(n894), .Z(n893) );
  OR2 C1854 ( .A(n900), .B(n895), .Z(n894) );
  OR2 C1853 ( .A(n901), .B(n902), .Z(n895) );
  IV I_25 ( .A(ENCODER_DATA_IN[49]), .Z(n896) );
  IV I_24 ( .A(ENCODER_DATA_IN[50]), .Z(n897) );
  IV I_23 ( .A(ENCODER_DATA_IN[51]), .Z(n898) );
  IV I_22 ( .A(ENCODER_DATA_IN[52]), .Z(n899) );
  IV I_21 ( .A(ENCODER_DATA_IN[53]), .Z(n900) );
  IV I_20 ( .A(ENCODER_DATA_IN[54]), .Z(n901) );
  IV I_19 ( .A(ENCODER_DATA_IN[55]), .Z(n902) );
  IV I_18 ( .A(n904), .Z(n903) );
  OR2 C1844 ( .A(ENCODER_DATA_IN[56]), .B(n905), .Z(n904) );
  OR2 C1843 ( .A(n911), .B(n906), .Z(n905) );
  OR2 C1842 ( .A(n912), .B(n907), .Z(n906) );
  OR2 C1841 ( .A(n913), .B(n908), .Z(n907) );
  OR2 C1840 ( .A(n914), .B(n909), .Z(n908) );
  OR2 C1839 ( .A(n915), .B(n910), .Z(n909) );
  OR2 C1838 ( .A(n916), .B(n917), .Z(n910) );
  IV I_17 ( .A(ENCODER_DATA_IN[57]), .Z(n911) );
  IV I_16 ( .A(ENCODER_DATA_IN[58]), .Z(n912) );
  IV I_15 ( .A(ENCODER_DATA_IN[59]), .Z(n913) );
  IV I_14 ( .A(ENCODER_DATA_IN[60]), .Z(n914) );
  IV I_13 ( .A(ENCODER_DATA_IN[61]), .Z(n915) );
  IV I_12 ( .A(ENCODER_DATA_IN[62]), .Z(n916) );
  IV I_11 ( .A(ENCODER_DATA_IN[63]), .Z(n917) );
  OR2 C1829 ( .A(U4_DATA1_0), .B(n920), .Z(n919) );
  OR2 C1828 ( .A(U4_DATA1_1), .B(n921), .Z(n920) );
  OR2 C1827 ( .A(U4_DATA1_2), .B(n922), .Z(n921) );
  OR2 C1826 ( .A(U4_DATA1_3), .B(n923), .Z(n922) );
  OR2 C1825 ( .A(U4_DATA1_4), .B(n924), .Z(n923) );
  OR2 C1824 ( .A(U4_DATA1_5), .B(n925), .Z(n924) );
  OR2 C1823 ( .A(U4_DATA1_6), .B(n926), .Z(n925) );
  OR2 C1822 ( .A(U4_DATA1_7), .B(U4_DATA1_8), .Z(n926) );
  OR2 C1817 ( .A(U4_DATA1_0), .B(n932), .Z(n931) );
  OR2 C1816 ( .A(U4_DATA1_1), .B(n933), .Z(n932) );
  OR2 C1815 ( .A(U4_DATA1_2), .B(n934), .Z(n933) );
  OR2 C1814 ( .A(U4_DATA1_3), .B(n935), .Z(n934) );
  OR2 C1813 ( .A(U4_DATA1_4), .B(n936), .Z(n935) );
  OR2 C1812 ( .A(U4_DATA1_5), .B(n937), .Z(n936) );
  OR2 C1811 ( .A(U4_DATA1_6), .B(n938), .Z(n937) );
  OR2 C1810 ( .A(n2460), .B(U4_DATA1_8), .Z(n938) );
  OR2 C1807 ( .A(U4_DATA1_0), .B(n941), .Z(n940) );
  OR2 C1806 ( .A(U4_DATA1_1), .B(n942), .Z(n941) );
  OR2 C1805 ( .A(U4_DATA1_2), .B(n943), .Z(n942) );
  OR2 C1804 ( .A(U4_DATA1_3), .B(n944), .Z(n943) );
  OR2 C1803 ( .A(U4_DATA1_4), .B(n945), .Z(n944) );
  OR2 C1802 ( .A(U4_DATA1_5), .B(n946), .Z(n945) );
  OR2 C1801 ( .A(U4_DATA1_6), .B(n947), .Z(n946) );
  OR2 C1800 ( .A(U4_DATA1_7), .B(n2412), .Z(n947) );
  OR2 C1797 ( .A(U4_DATA1_0), .B(n950), .Z(n949) );
  OR2 C1796 ( .A(U4_DATA1_1), .B(n951), .Z(n950) );
  OR2 C1795 ( .A(U4_DATA1_2), .B(n952), .Z(n951) );
  OR2 C1794 ( .A(U4_DATA1_3), .B(n953), .Z(n952) );
  OR2 C1793 ( .A(U4_DATA1_4), .B(n954), .Z(n953) );
  OR2 C1792 ( .A(U4_DATA1_5), .B(n955), .Z(n954) );
  OR2 C1791 ( .A(U4_DATA1_6), .B(n956), .Z(n955) );
  OR2 C1790 ( .A(n2460), .B(n2412), .Z(n956) );
  IV I_2 ( .A(n960), .Z(n959) );
  OR2 C1786 ( .A(ENCODER_CONTROL_IN[0]), .B(n961), .Z(n960) );
  OR2 C1785 ( .A(ENCODER_CONTROL_IN[1]), .B(n962), .Z(n961) );
  OR2 C1784 ( .A(ENCODER_CONTROL_IN[2]), .B(n963), .Z(n962) );
  OR2 C1783 ( .A(ENCODER_CONTROL_IN[3]), .B(n964), .Z(n963) );
  OR2 C1782 ( .A(ENCODER_CONTROL_IN[4]), .B(n965), .Z(n964) );
  OR2 C1781 ( .A(ENCODER_CONTROL_IN[5]), .B(n966), .Z(n965) );
  OR2 C1780 ( .A(ENCODER_CONTROL_IN[6]), .B(ENCODER_CONTROL_IN[7]), .Z(n966)
         );
  IV I_1 ( .A(RESET), .Z(n967) );
  IV I_0 ( .A(TEST_MODE), .Z(n968) );
  OR2 C1129 ( .A(n1444), .B(n1443), .Z(n1441) );
  OR2 C1128 ( .A(n1446), .B(n1445), .Z(n1442) );
  OR2 C1127 ( .A(n1447), .B(n[1743]), .Z(n1443) );
  OR2 C1126 ( .A(n1449), .B(n1448), .Z(n1444) );
  OR2 C1125 ( .A(n1451), .B(n1450), .Z(n1445) );
  OR2 C1124 ( .A(n1453), .B(n1452), .Z(n1446) );
  OR2 C1123 ( .A(n[1745]), .B(n[1744]), .Z(n1447) );
  OR2 C1122 ( .A(n[1747]), .B(n[1746]), .Z(n1448) );
  OR2 C1121 ( .A(n[1749]), .B(n[1748]), .Z(n1449) );
  OR2 C1120 ( .A(n[1751]), .B(n[1750]), .Z(n1450) );
  OR2 C1119 ( .A(n[1753]), .B(n[1752]), .Z(n1451) );
  OR2 C1118 ( .A(n[1755]), .B(n[1754]), .Z(n1452) );
  OR2 C1117 ( .A(n1454), .B(n[1756]), .Z(n1453) );
  OR2 C1113 ( .A(n1460), .B(n1459), .Z(n1457) );
  OR2 C1112 ( .A(n1462), .B(n1461), .Z(n1458) );
  OR2 C1111 ( .A(n1463), .B(n[1743]), .Z(n1459) );
  OR2 C1110 ( .A(n1465), .B(n1464), .Z(n1460) );
  OR2 C1109 ( .A(n1467), .B(n1466), .Z(n1461) );
  OR2 C1108 ( .A(n1469), .B(n1468), .Z(n1462) );
  OR2 C1107 ( .A(n[1745]), .B(n[1744]), .Z(n1463) );
  OR2 C1106 ( .A(n[1747]), .B(n[1746]), .Z(n1464) );
  OR2 C1105 ( .A(n[1749]), .B(n[1748]), .Z(n1465) );
  OR2 C1104 ( .A(n[1751]), .B(n[1750]), .Z(n1466) );
  OR2 C1103 ( .A(n[1753]), .B(n[1752]), .Z(n1467) );
  OR2 C1102 ( .A(n[1755]), .B(n[1754]), .Z(n1468) );
  OR2 C1101 ( .A(n[1757]), .B(n1470), .Z(n1469) );
  OR2 C1097 ( .A(n1476), .B(n1475), .Z(n1473) );
  OR2 C1096 ( .A(n1478), .B(n1477), .Z(n1474) );
  OR2 C1095 ( .A(n1479), .B(n[1743]), .Z(n1475) );
  OR2 C1094 ( .A(n1481), .B(n1480), .Z(n1476) );
  OR2 C1093 ( .A(n1483), .B(n1482), .Z(n1477) );
  OR2 C1092 ( .A(n1485), .B(n1484), .Z(n1478) );
  OR2 C1091 ( .A(n[1745]), .B(n[1744]), .Z(n1479) );
  OR2 C1090 ( .A(n[1747]), .B(n[1746]), .Z(n1480) );
  OR2 C1089 ( .A(n[1749]), .B(n[1748]), .Z(n1481) );
  OR2 C1088 ( .A(n[1751]), .B(n[1750]), .Z(n1482) );
  OR2 C1087 ( .A(n[1753]), .B(n[1752]), .Z(n1483) );
  OR2 C1086 ( .A(n1486), .B(n[1754]), .Z(n1484) );
  OR2 C1085 ( .A(n[1757]), .B(n[1756]), .Z(n1485) );
  OR2 C1081 ( .A(n1492), .B(n1491), .Z(n1489) );
  OR2 C1080 ( .A(n1494), .B(n1493), .Z(n1490) );
  OR2 C1079 ( .A(n1495), .B(n[1743]), .Z(n1491) );
  OR2 C1078 ( .A(n1497), .B(n1496), .Z(n1492) );
  OR2 C1077 ( .A(n1499), .B(n1498), .Z(n1493) );
  OR2 C1076 ( .A(n1501), .B(n1500), .Z(n1494) );
  OR2 C1075 ( .A(n[1745]), .B(n[1744]), .Z(n1495) );
  OR2 C1074 ( .A(n[1747]), .B(n[1746]), .Z(n1496) );
  OR2 C1073 ( .A(n[1749]), .B(n[1748]), .Z(n1497) );
  OR2 C1072 ( .A(n[1751]), .B(n[1750]), .Z(n1498) );
  OR2 C1071 ( .A(n[1753]), .B(n[1752]), .Z(n1499) );
  OR2 C1070 ( .A(n[1755]), .B(n1502), .Z(n1500) );
  OR2 C1069 ( .A(n[1757]), .B(n[1756]), .Z(n1501) );
  OR2 C1065 ( .A(n1508), .B(n1507), .Z(n1505) );
  OR2 C1064 ( .A(n1510), .B(n1509), .Z(n1506) );
  OR2 C1063 ( .A(n1511), .B(n[1743]), .Z(n1507) );
  OR2 C1062 ( .A(n1513), .B(n1512), .Z(n1508) );
  OR2 C1061 ( .A(n1515), .B(n1514), .Z(n1509) );
  OR2 C1060 ( .A(n1517), .B(n1516), .Z(n1510) );
  OR2 C1059 ( .A(n[1745]), .B(n[1744]), .Z(n1511) );
  OR2 C1058 ( .A(n[1747]), .B(n[1746]), .Z(n1512) );
  OR2 C1057 ( .A(n[1749]), .B(n[1748]), .Z(n1513) );
  OR2 C1056 ( .A(n[1751]), .B(n[1750]), .Z(n1514) );
  OR2 C1055 ( .A(n1518), .B(n[1752]), .Z(n1515) );
  OR2 C1054 ( .A(n[1755]), .B(n[1754]), .Z(n1516) );
  OR2 C1053 ( .A(n[1757]), .B(n[1756]), .Z(n1517) );
  OR2 C1049 ( .A(n1524), .B(n1523), .Z(n1521) );
  OR2 C1048 ( .A(n1526), .B(n1525), .Z(n1522) );
  OR2 C1047 ( .A(n1527), .B(n[1743]), .Z(n1523) );
  OR2 C1046 ( .A(n1529), .B(n1528), .Z(n1524) );
  OR2 C1045 ( .A(n1531), .B(n1530), .Z(n1525) );
  OR2 C1044 ( .A(n1533), .B(n1532), .Z(n1526) );
  OR2 C1043 ( .A(n[1745]), .B(n[1744]), .Z(n1527) );
  OR2 C1042 ( .A(n[1747]), .B(n[1746]), .Z(n1528) );
  OR2 C1041 ( .A(n[1749]), .B(n[1748]), .Z(n1529) );
  OR2 C1040 ( .A(n[1751]), .B(n[1750]), .Z(n1530) );
  OR2 C1039 ( .A(n[1753]), .B(n1534), .Z(n1531) );
  OR2 C1038 ( .A(n[1755]), .B(n[1754]), .Z(n1532) );
  OR2 C1037 ( .A(n[1757]), .B(n[1756]), .Z(n1533) );
  OR2 C1033 ( .A(n1540), .B(n1539), .Z(n1537) );
  OR2 C1032 ( .A(n1542), .B(n1541), .Z(n1538) );
  OR2 C1031 ( .A(n1543), .B(n[1743]), .Z(n1539) );
  OR2 C1030 ( .A(n1545), .B(n1544), .Z(n1540) );
  OR2 C1029 ( .A(n1547), .B(n1546), .Z(n1541) );
  OR2 C1028 ( .A(n1549), .B(n1548), .Z(n1542) );
  OR2 C1027 ( .A(n[1745]), .B(n[1744]), .Z(n1543) );
  OR2 C1026 ( .A(n[1747]), .B(n[1746]), .Z(n1544) );
  OR2 C1025 ( .A(n[1749]), .B(n[1748]), .Z(n1545) );
  OR2 C1024 ( .A(n1550), .B(n[1750]), .Z(n1546) );
  OR2 C1023 ( .A(n[1753]), .B(n[1752]), .Z(n1547) );
  OR2 C1022 ( .A(n[1755]), .B(n[1754]), .Z(n1548) );
  OR2 C1021 ( .A(n[1757]), .B(n[1756]), .Z(n1549) );
  OR2 C1017 ( .A(n1556), .B(n1555), .Z(n1553) );
  OR2 C1016 ( .A(n1558), .B(n1557), .Z(n1554) );
  OR2 C1015 ( .A(n1559), .B(n[1743]), .Z(n1555) );
  OR2 C1014 ( .A(n1561), .B(n1560), .Z(n1556) );
  OR2 C1013 ( .A(n1563), .B(n1562), .Z(n1557) );
  OR2 C1012 ( .A(n1565), .B(n1564), .Z(n1558) );
  OR2 C1011 ( .A(n[1745]), .B(n[1744]), .Z(n1559) );
  OR2 C1010 ( .A(n[1747]), .B(n[1746]), .Z(n1560) );
  OR2 C1009 ( .A(n[1749]), .B(n[1748]), .Z(n1561) );
  OR2 C1008 ( .A(n[1751]), .B(n1566), .Z(n1562) );
  OR2 C1007 ( .A(n[1753]), .B(n[1752]), .Z(n1563) );
  OR2 C1006 ( .A(n[1755]), .B(n[1754]), .Z(n1564) );
  OR2 C1005 ( .A(n[1757]), .B(n[1756]), .Z(n1565) );
  OR2 C1001 ( .A(n1572), .B(n1571), .Z(n1569) );
  OR2 C1000 ( .A(n1574), .B(n1573), .Z(n1570) );
  OR2 C999 ( .A(n1575), .B(n[1743]), .Z(n1571) );
  OR2 C998 ( .A(n1577), .B(n1576), .Z(n1572) );
  OR2 C997 ( .A(n1579), .B(n1578), .Z(n1573) );
  OR2 C996 ( .A(n1581), .B(n1580), .Z(n1574) );
  OR2 C995 ( .A(n[1745]), .B(n[1744]), .Z(n1575) );
  OR2 C994 ( .A(n[1747]), .B(n[1746]), .Z(n1576) );
  OR2 C993 ( .A(n1582), .B(n[1748]), .Z(n1577) );
  OR2 C992 ( .A(n[1751]), .B(n[1750]), .Z(n1578) );
  OR2 C991 ( .A(n[1753]), .B(n[1752]), .Z(n1579) );
  OR2 C990 ( .A(n[1755]), .B(n[1754]), .Z(n1580) );
  OR2 C989 ( .A(n[1757]), .B(n[1756]), .Z(n1581) );
  OR2 C985 ( .A(n1588), .B(n1587), .Z(n1585) );
  OR2 C984 ( .A(n1590), .B(n1589), .Z(n1586) );
  OR2 C983 ( .A(n1591), .B(n[1743]), .Z(n1587) );
  OR2 C982 ( .A(n1593), .B(n1592), .Z(n1588) );
  OR2 C981 ( .A(n1595), .B(n1594), .Z(n1589) );
  OR2 C980 ( .A(n1597), .B(n1596), .Z(n1590) );
  OR2 C979 ( .A(n[1745]), .B(n[1744]), .Z(n1591) );
  OR2 C978 ( .A(n[1747]), .B(n[1746]), .Z(n1592) );
  OR2 C977 ( .A(n[1749]), .B(n1598), .Z(n1593) );
  OR2 C976 ( .A(n[1751]), .B(n[1750]), .Z(n1594) );
  OR2 C975 ( .A(n[1753]), .B(n[1752]), .Z(n1595) );
  OR2 C974 ( .A(n[1755]), .B(n[1754]), .Z(n1596) );
  OR2 C973 ( .A(n[1757]), .B(n[1756]), .Z(n1597) );
  OR2 C969 ( .A(n1604), .B(n1603), .Z(n1601) );
  OR2 C968 ( .A(n1606), .B(n1605), .Z(n1602) );
  OR2 C967 ( .A(n1607), .B(n[1743]), .Z(n1603) );
  OR2 C966 ( .A(n1609), .B(n1608), .Z(n1604) );
  OR2 C965 ( .A(n1611), .B(n1610), .Z(n1605) );
  OR2 C964 ( .A(n1613), .B(n1612), .Z(n1606) );
  OR2 C963 ( .A(n[1745]), .B(n[1744]), .Z(n1607) );
  OR2 C962 ( .A(n1614), .B(n[1746]), .Z(n1608) );
  OR2 C961 ( .A(n[1749]), .B(n[1748]), .Z(n1609) );
  OR2 C960 ( .A(n[1751]), .B(n[1750]), .Z(n1610) );
  OR2 C959 ( .A(n[1753]), .B(n[1752]), .Z(n1611) );
  OR2 C958 ( .A(n[1755]), .B(n[1754]), .Z(n1612) );
  OR2 C957 ( .A(n[1757]), .B(n[1756]), .Z(n1613) );
  OR2 C953 ( .A(n1620), .B(n1619), .Z(n1617) );
  OR2 C952 ( .A(n1622), .B(n1621), .Z(n1618) );
  OR2 C951 ( .A(n1623), .B(n[1743]), .Z(n1619) );
  OR2 C950 ( .A(n1625), .B(n1624), .Z(n1620) );
  OR2 C949 ( .A(n1627), .B(n1626), .Z(n1621) );
  OR2 C948 ( .A(n1629), .B(n1628), .Z(n1622) );
  OR2 C947 ( .A(n[1745]), .B(n[1744]), .Z(n1623) );
  OR2 C946 ( .A(n[1747]), .B(n1630), .Z(n1624) );
  OR2 C945 ( .A(n[1749]), .B(n[1748]), .Z(n1625) );
  OR2 C944 ( .A(n[1751]), .B(n[1750]), .Z(n1626) );
  OR2 C943 ( .A(n[1753]), .B(n[1752]), .Z(n1627) );
  OR2 C942 ( .A(n[1755]), .B(n[1754]), .Z(n1628) );
  OR2 C941 ( .A(n[1757]), .B(n[1756]), .Z(n1629) );
  OR2 C937 ( .A(n1636), .B(n1635), .Z(n1633) );
  OR2 C936 ( .A(n1638), .B(n1637), .Z(n1634) );
  OR2 C935 ( .A(n1639), .B(n[1743]), .Z(n1635) );
  OR2 C934 ( .A(n1641), .B(n1640), .Z(n1636) );
  OR2 C933 ( .A(n1643), .B(n1642), .Z(n1637) );
  OR2 C932 ( .A(n1645), .B(n1644), .Z(n1638) );
  OR2 C931 ( .A(n1646), .B(n[1744]), .Z(n1639) );
  OR2 C930 ( .A(n[1747]), .B(n[1746]), .Z(n1640) );
  OR2 C929 ( .A(n[1749]), .B(n[1748]), .Z(n1641) );
  OR2 C928 ( .A(n[1751]), .B(n[1750]), .Z(n1642) );
  OR2 C927 ( .A(n[1753]), .B(n[1752]), .Z(n1643) );
  OR2 C926 ( .A(n[1755]), .B(n[1754]), .Z(n1644) );
  OR2 C925 ( .A(n[1757]), .B(n[1756]), .Z(n1645) );
  OR2 C921 ( .A(n1652), .B(n1651), .Z(n1649) );
  OR2 C920 ( .A(n1654), .B(n1653), .Z(n1650) );
  OR2 C919 ( .A(n1655), .B(n[1743]), .Z(n1651) );
  OR2 C918 ( .A(n1657), .B(n1656), .Z(n1652) );
  OR2 C917 ( .A(n1659), .B(n1658), .Z(n1653) );
  OR2 C916 ( .A(n1661), .B(n1660), .Z(n1654) );
  OR2 C915 ( .A(n[1745]), .B(n1662), .Z(n1655) );
  OR2 C914 ( .A(n[1747]), .B(n[1746]), .Z(n1656) );
  OR2 C913 ( .A(n[1749]), .B(n[1748]), .Z(n1657) );
  OR2 C912 ( .A(n[1751]), .B(n[1750]), .Z(n1658) );
  OR2 C911 ( .A(n[1753]), .B(n[1752]), .Z(n1659) );
  OR2 C910 ( .A(n[1755]), .B(n[1754]), .Z(n1660) );
  OR2 C909 ( .A(n[1757]), .B(n[1756]), .Z(n1661) );
  OR2 C905 ( .A(n1668), .B(n1667), .Z(n1665) );
  OR2 C904 ( .A(n1670), .B(n1669), .Z(n1666) );
  OR2 C903 ( .A(n1671), .B(n1678), .Z(n1667) );
  OR2 C902 ( .A(n1673), .B(n1672), .Z(n1668) );
  OR2 C901 ( .A(n1675), .B(n1674), .Z(n1669) );
  OR2 C900 ( .A(n1677), .B(n1676), .Z(n1670) );
  OR2 C899 ( .A(n[1745]), .B(n[1744]), .Z(n1671) );
  OR2 C898 ( .A(n[1747]), .B(n[1746]), .Z(n1672) );
  OR2 C897 ( .A(n[1749]), .B(n[1748]), .Z(n1673) );
  OR2 C896 ( .A(n[1751]), .B(n[1750]), .Z(n1674) );
  OR2 C895 ( .A(n[1753]), .B(n[1752]), .Z(n1675) );
  OR2 C894 ( .A(n[1755]), .B(n[1754]), .Z(n1676) );
  OR2 C893 ( .A(n[1757]), .B(n[1756]), .Z(n1677) );
  FD1 drs1_reg ( .D(DATA_PAT_SEL), .CP(CLK), .Q(n6) );
  FD1 drs2_reg ( .D(n6), .CP(CLK), .Q(n1971) );
  FD1 drs1_reg1 ( .D(TEST_MODE), .CP(CLK), .Q(n3) );
  FD1 drs2_reg1 ( .D(n3), .CP(CLK), .Q(n1970) );
  FD1 test_counter_reg_0_ ( .D(U6_Z_0), .CP(CLK), .Q(U4_DATA1_0) );
  FD1 test_counter_reg_1_ ( .D(U6_Z_1), .CP(CLK), .Q(U4_DATA1_1) );
  FD1 test_counter_reg_2_ ( .D(U6_Z_2), .CP(CLK), .Q(U4_DATA1_2) );
  FD1 test_counter_reg_3_ ( .D(U6_Z_3), .CP(CLK), .Q(U4_DATA1_3) );
  FD1 test_counter_reg_4_ ( .D(U6_Z_4), .CP(CLK), .Q(U4_DATA1_4) );
  FD1 test_counter_reg_5_ ( .D(U6_Z_5), .CP(CLK), .Q(U4_DATA1_5) );
  FD1 test_counter_reg_6_ ( .D(U6_Z_6), .CP(CLK), .Q(U4_DATA1_6) );
  FD1 test_counter_reg_7_ ( .D(U6_Z_7), .CP(CLK), .Q(U4_DATA1_7) );
  FD1 test_counter_reg_8_ ( .D(U6_Z_8), .CP(CLK), .Q(U4_DATA1_8) );
  FD1 data_prev_reg_9_ ( .D(U5_Z_9), .CP(CLK), .Q(U7_DATA1_9) );
  FD1 data_prev_reg_3_ ( .D(U5_Z_3), .CP(CLK), .Q(U7_DATA1_3) );
  FD1 data_prev_reg_42_ ( .D(U5_Z_42), .CP(CLK), .Q(U7_DATA1_42) );
  FD1 data_prev_reg_36_ ( .D(U5_Z_36), .CP(CLK), .Q(U7_DATA1_36) );
  FD1 data_prev_reg_30_ ( .D(U5_Z_30), .CP(CLK), .Q(U7_DATA1_30) );
  FD1 data_prev_reg_5_ ( .D(U5_Z_5), .CP(CLK), .Q(U7_DATA1_5) );
  FD1 data_prev_reg_57_ ( .D(U5_Z_57), .CP(CLK), .Q(U7_DATA1_57) );
  FD1 data_prev_reg_51_ ( .D(U5_Z_51), .CP(CLK), .Q(U7_DATA1_51) );
  FD1 data_prev_reg_45_ ( .D(U5_Z_45), .CP(CLK), .Q(U7_DATA1_45) );
  FD1 data_prev_reg_39_ ( .D(U5_Z_39), .CP(CLK), .Q(U7_DATA1_39) );
  FD1 data_prev_reg_33_ ( .D(U5_Z_33), .CP(CLK), .Q(U7_DATA1_33) );
  FD1 data_prev_reg_8_ ( .D(U5_Z_8), .CP(CLK), .Q(U7_DATA1_8) );
  FD1 data_prev_reg_2_ ( .D(U5_Z_2), .CP(CLK), .Q(U7_DATA1_2) );
  FD1 data_prev_reg_41_ ( .D(U5_Z_41), .CP(CLK), .Q(U7_DATA1_41) );
  FD1 data_prev_reg_35_ ( .D(U5_Z_35), .CP(CLK), .Q(U7_DATA1_35) );
  FD1 data_prev_reg_29_ ( .D(U5_Z_29), .CP(CLK), .Q(U7_DATA1_29) );
  FD1 data_prev_reg_4_ ( .D(U5_Z_4), .CP(CLK), .Q(U7_DATA1_4) );
  FD1 data_prev_reg_43_ ( .D(U5_Z_43), .CP(CLK), .Q(U7_DATA1_43) );
  FD1 data_prev_reg_37_ ( .D(U5_Z_37), .CP(CLK), .Q(U7_DATA1_37) );
  FD1 data_prev_reg_31_ ( .D(U5_Z_31), .CP(CLK), .Q(U7_DATA1_31) );
  FD1 data_prev_reg_6_ ( .D(U5_Z_6), .CP(CLK), .Q(U7_DATA1_6) );
  FD1 data_prev_reg_0_ ( .D(U5_Z_0), .CP(CLK), .Q(U7_DATA1_0) );
  FD1 data_prev_reg_52_ ( .D(U5_Z_52), .CP(CLK), .Q(U7_DATA1_52) );
  FD1 data_prev_reg_27_ ( .D(U5_Z_27), .CP(CLK), .Q(U7_DATA1_27) );
  FD1 data_prev_reg_46_ ( .D(U5_Z_46), .CP(CLK), .Q(U7_DATA1_46) );
  FD1 data_prev_reg_21_ ( .D(U5_Z_21), .CP(CLK), .Q(U7_DATA1_21) );
  FD1 data_prev_reg_40_ ( .D(U5_Z_40), .CP(CLK), .Q(U7_DATA1_40) );
  FD1 data_prev_reg_15_ ( .D(U5_Z_15), .CP(CLK), .Q(U7_DATA1_15) );
  FD1 data_prev_reg_54_ ( .D(U5_Z_54), .CP(CLK), .Q(U7_DATA1_54) );
  FD1 data_prev_reg_34_ ( .D(U5_Z_34), .CP(CLK), .Q(U7_DATA1_34) );
  FD1 data_prev_reg_48_ ( .D(U5_Z_48), .CP(CLK), .Q(U7_DATA1_48) );
  FD1 data_prev_reg_23_ ( .D(U5_Z_23), .CP(CLK), .Q(U7_DATA1_23) );
  FD1 data_prev_reg_17_ ( .D(U5_Z_17), .CP(CLK), .Q(U7_DATA1_17) );
  FD1 data_prev_reg_11_ ( .D(U5_Z_11), .CP(CLK), .Q(U7_DATA1_11) );
  FD1 data_prev_reg_56_ ( .D(U5_Z_56), .CP(CLK), .Q(U7_DATA1_56) );
  FD1 data_prev_reg_50_ ( .D(U5_Z_50), .CP(CLK), .Q(U7_DATA1_50) );
  FD1 data_prev_reg_25_ ( .D(U5_Z_25), .CP(CLK), .Q(U7_DATA1_25) );
  FD1 data_prev_reg_44_ ( .D(U5_Z_44), .CP(CLK), .Q(U7_DATA1_44) );
  FD1 data_prev_reg_19_ ( .D(U5_Z_19), .CP(CLK), .Q(U7_DATA1_19) );
  FD1 data_prev_reg_38_ ( .D(U5_Z_38), .CP(CLK), .Q(U7_DATA1_38) );
  FD1 data_prev_reg_13_ ( .D(U5_Z_13), .CP(CLK), .Q(U7_DATA1_13) );
  FD1 data_prev_reg_32_ ( .D(U5_Z_32), .CP(CLK), .Q(U7_DATA1_32) );
  FD1 data_prev_reg_26_ ( .D(U5_Z_26), .CP(CLK), .Q(U7_DATA1_26) );
  FD1 data_prev_reg_20_ ( .D(U5_Z_20), .CP(CLK), .Q(U7_DATA1_20) );
  FD1 data_prev_reg_14_ ( .D(U5_Z_14), .CP(CLK), .Q(U7_DATA1_14) );
  FD1 data_prev_reg_7_ ( .D(U5_Z_7), .CP(CLK), .Q(U7_DATA1_7) );
  FD1 data_prev_reg_1_ ( .D(U5_Z_1), .CP(CLK), .Q(U7_DATA1_1) );
  FD1 data_prev_reg_53_ ( .D(U5_Z_53), .CP(CLK), .Q(U7_DATA1_53) );
  FD1 data_prev_reg_28_ ( .D(U5_Z_28), .CP(CLK), .Q(U7_DATA1_28) );
  FD1 data_prev_reg_47_ ( .D(U5_Z_47), .CP(CLK), .Q(U7_DATA1_47) );
  FD1 data_prev_reg_22_ ( .D(U5_Z_22), .CP(CLK), .Q(U7_DATA1_22) );
  FD1 data_prev_reg_16_ ( .D(U5_Z_16), .CP(CLK), .Q(U7_DATA1_16) );
  FD1 data_prev_reg_10_ ( .D(U5_Z_10), .CP(CLK), .Q(U7_DATA1_10) );
  FD1 data_prev_reg_55_ ( .D(U5_Z_55), .CP(CLK), .Q(U7_DATA1_55) );
  FD1 data_prev_reg_49_ ( .D(U5_Z_49), .CP(CLK), .Q(U7_DATA1_49) );
  FD1 data_prev_reg_24_ ( .D(U5_Z_24), .CP(CLK), .Q(U7_DATA1_24) );
  FD1 data_prev_reg_18_ ( .D(U5_Z_18), .CP(CLK), .Q(U7_DATA1_18) );
  FD1 data_prev_reg_12_ ( .D(U5_Z_12), .CP(CLK), .Q(U7_DATA1_12) );
  IV U196 ( .A(DATA_VALID), .Z(n2474) );
  IV U197 ( .A(n1759), .Z(n2475) );
  IV U198 ( .A(n1760), .Z(n2476) );
  IV U199 ( .A(n2586), .Z(n2477) );
  IV U200 ( .A(n2587), .Z(n2478) );
  IV U201 ( .A(n2590), .Z(n2479) );
  IV U202 ( .A(n2588), .Z(n2480) );
  IV U203 ( .A(n2592), .Z(n2481) );
  IV U204 ( .A(n1772), .Z(n2482) );
  IV U205 ( .A(n2593), .Z(n2483) );
  IV U206 ( .A(n2595), .Z(n2484) );
  IV U207 ( .A(n2597), .Z(n2485) );
  IV U208 ( .A(n1944), .Z(n2486) );
  IV U209 ( .A(n1770), .Z(n2487) );
  IV U210 ( .A(n1768), .Z(n2488) );
  OR2 U214 ( .A(n1535), .B(n2560), .Z(n328) );
  OR2 U215 ( .A(n2561), .B(n2562), .Z(n327) );
  OR2 U216 ( .A(n1615), .B(n2563), .Z(n2562) );
  OR2 U217 ( .A(n1663), .B(n1631), .Z(n2561) );
  OR2 U218 ( .A(n2564), .B(n2565), .Z(n326) );
  OR2 U219 ( .A(n1519), .B(n1471), .Z(n2565) );
  OR2 U220 ( .A(n2566), .B(n2567), .Z(n325) );
  OR2 U221 ( .A(n1551), .B(n2568), .Z(n2567) );
  OR2 U222 ( .A(n1663), .B(n1647), .Z(n2566) );
  OR2 U223 ( .A(n2569), .B(n2564), .Z(n324) );
  OR2 U224 ( .A(n2570), .B(n2571), .Z(n323) );
  OR2 U225 ( .A(n1567), .B(n2572), .Z(n2571) );
  OR2 U226 ( .A(n1647), .B(n1583), .Z(n2570) );
  OR2 U227 ( .A(n2564), .B(n2573), .Z(n322) );
  OR2 U228 ( .A(n1519), .B(n1487), .Z(n2573) );
  OR2 U229 ( .A(n2574), .B(n2575), .Z(n321) );
  OR2 U230 ( .A(n1583), .B(n2572), .Z(n2575) );
  OR2 U231 ( .A(n1631), .B(n1599), .Z(n2574) );
  OR2 U232 ( .A(n2564), .B(n2576), .Z(n320) );
  OR2 U233 ( .A(n1503), .B(n1471), .Z(n2576) );
  OR2 U234 ( .A(U33_CONTROL5), .B(n1439), .Z(n2564) );
  OR2 U235 ( .A(n2577), .B(n2578), .Z(n319) );
  OR2 U236 ( .A(n1519), .B(n2579), .Z(n2578) );
  OR2 U237 ( .A(n1615), .B(n1583), .Z(n2577) );
  OR2 U238 ( .A(n1503), .B(n2560), .Z(n318) );
  OR2 U239 ( .A(n1487), .B(U34_CONTROL2), .Z(n316) );
  OR2 U240 ( .A(n2580), .B(n2581), .Z(n314) );
  OR2 U241 ( .A(n1519), .B(n2569), .Z(n2581) );
  OR2 U242 ( .A(n1551), .B(n1535), .Z(n2580) );
  OR2 U243 ( .A(n1519), .B(n284), .Z(n306) );
  OR2 U244 ( .A(n2572), .B(n2582), .Z(n297) );
  OR2 U245 ( .A(n1519), .B(n2563), .Z(n2582) );
  OR2 U246 ( .A(n1535), .B(n1663), .Z(n2572) );
  OR2 U247 ( .A(n1455), .B(n287), .Z(n284) );
  AN2 U248 ( .A(n2583), .B(n2584), .Z(n[1757]) );
  AN2 U249 ( .A(n2475), .B(n2476), .Z(n2584) );
  AN2 U250 ( .A(n1758), .B(n2477), .Z(n2583) );
  AN2 U251 ( .A(n2585), .B(n1759), .Z(n[1756]) );
  AN2 U252 ( .A(n2477), .B(n2476), .Z(n2585) );
  AN2 U253 ( .A(n1760), .B(n2477), .Z(n[1755]) );
  OR2 U254 ( .A(n1761), .B(n2587), .Z(n2586) );
  AN2 U255 ( .A(n1761), .B(n2478), .Z(n[1754]) );
  OR2 U256 ( .A(n2588), .B(n2589), .Z(n2587) );
  OR2 U257 ( .A(n1763), .B(n1762), .Z(n2589) );
  AN2 U258 ( .A(n2479), .B(n1762), .Z(n[1753]) );
  OR2 U259 ( .A(n2588), .B(n1763), .Z(n2590) );
  AN2 U260 ( .A(n1763), .B(n2480), .Z(n[1752]) );
  OR2 U261 ( .A(n1764), .B(n2591), .Z(n2588) );
  AN2 U262 ( .A(n1764), .B(U3_n725), .Z(n[1751]) );
  AN2 U263 ( .A(n2481), .B(n1765), .Z(n[1750]) );
  OR2 U264 ( .A(n2593), .B(n1766), .Z(n2592) );
  AN2 U265 ( .A(n1766), .B(n2483), .Z(n[1749]) );
  AN2 U266 ( .A(n2594), .B(n1767), .Z(n[1748]) );
  AN2 U267 ( .A(n2484), .B(n2488), .Z(n2594) );
  AN2 U268 ( .A(n1768), .B(n2484), .Z(n[1747]) );
  AN2 U269 ( .A(n2596), .B(n1769), .Z(n[1746]) );
  AN2 U270 ( .A(n2485), .B(n2487), .Z(n2596) );
  AN2 U271 ( .A(n1770), .B(n2485), .Z(n[1745]) );
  AN2 U272 ( .A(n2598), .B(n1771), .Z(n[1744]) );
  AN2 U273 ( .A(n2482), .B(n2486), .Z(n2598) );
  AN2 U274 ( .A(n1772), .B(n2486), .Z(n[1743]) );
  OR2 U275 ( .A(n1665), .B(n1666), .Z(n1664) );
  OR2 U276 ( .A(n1649), .B(n1650), .Z(n1648) );
  OR2 U277 ( .A(n1633), .B(n1634), .Z(n1632) );
  OR2 U278 ( .A(n1617), .B(n1618), .Z(n1616) );
  OR2 U279 ( .A(n1601), .B(n1602), .Z(n1600) );
  OR2 U280 ( .A(n1585), .B(n1586), .Z(n1584) );
  OR2 U281 ( .A(n1569), .B(n1570), .Z(n1568) );
  OR2 U282 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR2 U283 ( .A(n1537), .B(n1538), .Z(n1536) );
  OR2 U284 ( .A(n1521), .B(n1522), .Z(n1520) );
  OR2 U285 ( .A(n1505), .B(n1506), .Z(n1504) );
  OR2 U286 ( .A(n1489), .B(n1490), .Z(n1488) );
  OR2 U287 ( .A(n1473), .B(n1474), .Z(n1472) );
  OR2 U288 ( .A(n1457), .B(n1458), .Z(n1456) );
  OR2 U289 ( .A(n1441), .B(n1442), .Z(n1440) );
  AN2 U1561 ( .A(n1046), .B(n967), .Z(n2661) );
  OR2 U1590 ( .A(n2474), .B(RESET), .Z(n3749) );
  OR2 U1593 ( .A(n3773), .B(n3774), .Z(U34_Z_2) );
  OR2 U1594 ( .A(n3775), .B(n3776), .Z(n3774) );
  AN2 U1595 ( .A(ENCODER_DATA_IN[14]), .B(U34_CONTROL2), .Z(n3776) );
  AN2 U1596 ( .A(U34_DATA1_2), .B(U34_CONTROL1), .Z(n3775) );
  AN2 U1597 ( .A(ENCODER_DATA_IN[6]), .B(n308), .Z(n3773) );
  OR2 U1598 ( .A(n3777), .B(n3778), .Z(U34_Z_1) );
  OR2 U1599 ( .A(n3779), .B(n3780), .Z(n3778) );
  AN2 U1600 ( .A(ENCODER_DATA_IN[13]), .B(U34_CONTROL2), .Z(n3780) );
  AN2 U1601 ( .A(U34_DATA1_1), .B(U34_CONTROL1), .Z(n3779) );
  AN2 U1602 ( .A(ENCODER_DATA_IN[5]), .B(n308), .Z(n3777) );
  OR2 U1603 ( .A(n3781), .B(n3782), .Z(U34_Z_0) );
  OR2 U1604 ( .A(n3783), .B(n3784), .Z(n3782) );
  AN2 U1605 ( .A(ENCODER_DATA_IN[8]), .B(U34_CONTROL2), .Z(n3784) );
  AN2 U1606 ( .A(U34_DATA1_0), .B(U34_CONTROL1), .Z(n3783) );
  AN2 U1607 ( .A(ENCODER_DATA_IN[0]), .B(n308), .Z(n3781) );
  OR2 U1608 ( .A(n3785), .B(n3786), .Z(U34_DATA1_2) );
  OR2 U1609 ( .A(n3787), .B(n3786), .Z(U34_DATA1_1) );
  OR2 U1610 ( .A(n1931), .B(n1930), .Z(n3786) );
  OR2 U1611 ( .A(n3785), .B(n3787), .Z(U34_DATA1_0) );
  OR2 U1612 ( .A(n1933), .B(n1932), .Z(n3787) );
  OR2 U1613 ( .A(n1935), .B(n1934), .Z(n3785) );
  OR2 U1614 ( .A(n3788), .B(n3789), .Z(U33_Z_3) );
  OR2 U1615 ( .A(n3790), .B(n3791), .Z(n3789) );
  AN2 U1616 ( .A(ENCODER_DATA_IN[4]), .B(n308), .Z(n3791) );
  AN2 U1617 ( .A(ENCODER_DATA_IN[12]), .B(U34_CONTROL2), .Z(n3790) );
  OR2 U1618 ( .A(U33_CONTROL5), .B(n3792), .Z(n3788) );
  AN2 U1619 ( .A(U33_DATA1_3), .B(U34_CONTROL1), .Z(n3792) );
  OR2 U1620 ( .A(n3793), .B(n3794), .Z(U33_Z_2) );
  OR2 U1621 ( .A(n3795), .B(n3796), .Z(n3794) );
  AN2 U1622 ( .A(ENCODER_DATA_IN[3]), .B(n308), .Z(n3796) );
  AN2 U1623 ( .A(ENCODER_DATA_IN[11]), .B(U34_CONTROL2), .Z(n3795) );
  OR2 U1624 ( .A(U33_CONTROL5), .B(n3797), .Z(n3793) );
  AN2 U1625 ( .A(U33_DATA1_2), .B(U34_CONTROL1), .Z(n3797) );
  OR2 U1626 ( .A(n3798), .B(n3799), .Z(U33_Z_1) );
  OR2 U1627 ( .A(n3800), .B(n3801), .Z(n3799) );
  AN2 U1628 ( .A(ENCODER_DATA_IN[2]), .B(n308), .Z(n3801) );
  AN2 U1629 ( .A(ENCODER_DATA_IN[10]), .B(U34_CONTROL2), .Z(n3800) );
  OR2 U1630 ( .A(U33_CONTROL5), .B(n3802), .Z(n3798) );
  AN2 U1631 ( .A(U33_DATA1_1), .B(U34_CONTROL1), .Z(n3802) );
  OR2 U1632 ( .A(n3803), .B(n3804), .Z(U33_Z_0) );
  OR2 U1633 ( .A(n3805), .B(n3806), .Z(n3804) );
  AN2 U1634 ( .A(ENCODER_DATA_IN[1]), .B(n308), .Z(n3806) );
  AN2 U1635 ( .A(ENCODER_DATA_IN[9]), .B(U34_CONTROL2), .Z(n3805) );
  OR2 U1636 ( .A(U33_CONTROL5), .B(n3807), .Z(n3803) );
  AN2 U1637 ( .A(U33_DATA1_0), .B(U34_CONTROL1), .Z(n3807) );
  OR2 U1638 ( .A(n3808), .B(n3809), .Z(U33_DATA1_3) );
  OR2 U1639 ( .A(n1934), .B(n1932), .Z(n3808) );
  OR2 U1640 ( .A(n3810), .B(n3809), .Z(U33_DATA1_2) );
  OR2 U1641 ( .A(n1930), .B(n3811), .Z(n3809) );
  AN2 U1642 ( .A(n3812), .B(n720), .Z(n1930) );
  OR2 U1643 ( .A(n1935), .B(n1933), .Z(n3810) );
  OR2 U1644 ( .A(n3813), .B(n3814), .Z(U33_DATA1_1) );
  OR2 U1645 ( .A(n1934), .B(n1933), .Z(n3813) );
  AN2 U1646 ( .A(n542), .B(n3815), .Z(n1933) );
  AN2 U1647 ( .A(n3816), .B(n478), .Z(n1934) );
  OR2 U1648 ( .A(n3817), .B(n3814), .Z(U33_DATA1_0) );
  OR2 U1649 ( .A(n1931), .B(n3811), .Z(n3814) );
  OR2 U1650 ( .A(n1929), .B(n1943), .Z(n3811) );
  IV U1651 ( .A(n3818), .Z(n1943) );
  OR2 U1652 ( .A(n3819), .B(n3820), .Z(n3818) );
  OR2 U1653 ( .A(n3821), .B(n3822), .Z(n3820) );
  OR2 U1654 ( .A(n377), .B(n376), .Z(n3822) );
  OR2 U1655 ( .A(n478), .B(n418), .Z(n3821) );
  OR2 U1656 ( .A(n3823), .B(n3824), .Z(n3819) );
  OR2 U1657 ( .A(n600), .B(n542), .Z(n3824) );
  OR2 U1658 ( .A(n662), .B(n3825), .Z(n3823) );
  OR2 U1659 ( .A(n770), .B(n720), .Z(n3825) );
  AN2 U1660 ( .A(n770), .B(n3826), .Z(n1929) );
  AN2 U1661 ( .A(n3812), .B(n721), .Z(n3826) );
  AN2 U1662 ( .A(n3827), .B(n663), .Z(n3812) );
  AN2 U1663 ( .A(n662), .B(n3827), .Z(n1931) );
  AN2 U1664 ( .A(n601), .B(n3828), .Z(n3827) );
  OR2 U1665 ( .A(n1935), .B(n1932), .Z(n3817) );
  AN2 U1666 ( .A(n3828), .B(n600), .Z(n1932) );
  AN2 U1667 ( .A(n543), .B(n3815), .Z(n3828) );
  AN2 U1668 ( .A(n3816), .B(n479), .Z(n3815) );
  AN2 U1669 ( .A(n419), .B(n3829), .Z(n3816) );
  AN2 U1670 ( .A(n418), .B(n3829), .Z(n1935) );
  AN2 U1671 ( .A(ENCODER_CONTROL_IN[0]), .B(n378), .Z(n3829) );
  OR2 U1672 ( .A(n3830), .B(n3831), .Z(U32_Z_0) );
  OR2 U1673 ( .A(n3832), .B(n3833), .Z(n3831) );
  AN2 U1674 ( .A(ENCODER_DATA_IN[15]), .B(U34_CONTROL2), .Z(n3833) );
  AN2 U1675 ( .A(U32_DATA1_0), .B(U32_CONTROL1), .Z(n3832) );
  AN2 U1676 ( .A(n308), .B(ENCODER_DATA_IN[7]), .Z(n3830) );
  OR2 U1677 ( .A(n3834), .B(n3835), .Z(U32_DATA1_0) );
  OR2 U1678 ( .A(n3836), .B(n3837), .Z(U31_Z_3) );
  OR2 U1679 ( .A(n3838), .B(n3839), .Z(n3837) );
  AN2 U1680 ( .A(ENCODER_DATA_IN[11]), .B(n305), .Z(n3839) );
  AN2 U1681 ( .A(ENCODER_DATA_IN[19]), .B(U34_CONTROL2), .Z(n3838) );
  OR2 U1682 ( .A(U33_CONTROL5), .B(n3840), .Z(n3836) );
  AN2 U1683 ( .A(U31_DATA1_3), .B(U32_CONTROL1), .Z(n3840) );
  OR2 U1684 ( .A(n3841), .B(n3842), .Z(U31_Z_2) );
  OR2 U1685 ( .A(n3843), .B(n3844), .Z(n3842) );
  AN2 U1686 ( .A(ENCODER_DATA_IN[10]), .B(n305), .Z(n3844) );
  AN2 U1687 ( .A(ENCODER_DATA_IN[18]), .B(U34_CONTROL2), .Z(n3843) );
  OR2 U1688 ( .A(U33_CONTROL5), .B(n3845), .Z(n3841) );
  AN2 U1689 ( .A(U31_DATA1_2), .B(U32_CONTROL1), .Z(n3845) );
  OR2 U1690 ( .A(n3846), .B(n3847), .Z(U31_Z_1) );
  OR2 U1691 ( .A(n3848), .B(n3849), .Z(n3847) );
  AN2 U1692 ( .A(ENCODER_DATA_IN[9]), .B(n305), .Z(n3849) );
  AN2 U1693 ( .A(ENCODER_DATA_IN[17]), .B(U34_CONTROL2), .Z(n3848) );
  OR2 U1694 ( .A(U33_CONTROL5), .B(n3850), .Z(n3846) );
  AN2 U1695 ( .A(U31_DATA1_1), .B(U32_CONTROL1), .Z(n3850) );
  OR2 U1696 ( .A(n3851), .B(n3852), .Z(U31_Z_0) );
  OR2 U1697 ( .A(n3853), .B(n3854), .Z(n3852) );
  AN2 U1698 ( .A(ENCODER_DATA_IN[8]), .B(n305), .Z(n3854) );
  AN2 U1699 ( .A(ENCODER_DATA_IN[16]), .B(U34_CONTROL2), .Z(n3853) );
  OR2 U1700 ( .A(U33_CONTROL5), .B(n3855), .Z(n3851) );
  AN2 U1701 ( .A(U31_DATA1_0), .B(U32_CONTROL1), .Z(n3855) );
  OR2 U1702 ( .A(n3856), .B(n3857), .Z(U31_DATA1_3) );
  OR2 U1703 ( .A(n1919), .B(n1917), .Z(n3856) );
  OR2 U1704 ( .A(n3858), .B(n3857), .Z(U31_DATA1_2) );
  OR2 U1705 ( .A(n1915), .B(n3859), .Z(n3857) );
  OR2 U1706 ( .A(n1920), .B(n1918), .Z(n3858) );
  OR2 U1707 ( .A(n3860), .B(n3861), .Z(U31_DATA1_1) );
  OR2 U1708 ( .A(n1919), .B(n1918), .Z(n3860) );
  OR2 U1709 ( .A(n3862), .B(n3861), .Z(U31_DATA1_0) );
  OR2 U1710 ( .A(n1916), .B(n3859), .Z(n3861) );
  OR2 U1711 ( .A(n1914), .B(n1928), .Z(n3859) );
  IV U1712 ( .A(n3863), .Z(n1928) );
  OR2 U1713 ( .A(n3864), .B(n3865), .Z(n3863) );
  OR2 U1714 ( .A(n3866), .B(n3867), .Z(n3865) );
  OR2 U1715 ( .A(n384), .B(n383), .Z(n3867) );
  OR2 U1716 ( .A(n494), .B(n432), .Z(n3866) );
  OR2 U1717 ( .A(n3868), .B(n3869), .Z(n3864) );
  OR2 U1718 ( .A(n615), .B(n557), .Z(n3869) );
  OR2 U1719 ( .A(n677), .B(n3870), .Z(n3868) );
  OR2 U1720 ( .A(n787), .B(n733), .Z(n3870) );
  AN2 U1721 ( .A(n787), .B(n3871), .Z(n1914) );
  AN2 U1722 ( .A(n3872), .B(n734), .Z(n3871) );
  OR2 U1723 ( .A(n1920), .B(n1917), .Z(n3862) );
  OR2 U1724 ( .A(n3873), .B(n3874), .Z(U30_Z_1) );
  OR2 U1725 ( .A(n3875), .B(n3876), .Z(n3874) );
  AN2 U1726 ( .A(ENCODER_DATA_IN[21]), .B(U34_CONTROL2), .Z(n3876) );
  AN2 U1727 ( .A(U30_DATA1_1), .B(U32_CONTROL1), .Z(n3875) );
  AN2 U1728 ( .A(n305), .B(ENCODER_DATA_IN[13]), .Z(n3873) );
  OR2 U1729 ( .A(n3877), .B(n3878), .Z(U30_Z_0) );
  OR2 U1730 ( .A(n3879), .B(n3880), .Z(n3878) );
  AN2 U1731 ( .A(ENCODER_DATA_IN[20]), .B(U34_CONTROL2), .Z(n3880) );
  AN2 U1732 ( .A(U30_DATA1_0), .B(U32_CONTROL1), .Z(n3879) );
  AN2 U1733 ( .A(n305), .B(ENCODER_DATA_IN[12]), .Z(n3877) );
  OR2 U1734 ( .A(n3834), .B(n3881), .Z(U30_DATA1_1) );
  OR2 U1735 ( .A(n1920), .B(n1919), .Z(n3834) );
  AN2 U1736 ( .A(n3882), .B(n494), .Z(n1919) );
  AN2 U1737 ( .A(n432), .B(n3883), .Z(n1920) );
  OR2 U1738 ( .A(n3835), .B(n3881), .Z(U30_DATA1_0) );
  OR2 U1739 ( .A(n1916), .B(n1915), .Z(n3881) );
  AN2 U1740 ( .A(n3872), .B(n733), .Z(n1915) );
  AN2 U1741 ( .A(n3884), .B(n678), .Z(n3872) );
  AN2 U1742 ( .A(n677), .B(n3884), .Z(n1916) );
  AN2 U1743 ( .A(n616), .B(n3885), .Z(n3884) );
  OR2 U1744 ( .A(n1918), .B(n1917), .Z(n3835) );
  AN2 U1745 ( .A(n3885), .B(n615), .Z(n1917) );
  AN2 U1746 ( .A(n558), .B(n3886), .Z(n3885) );
  AN2 U1747 ( .A(n557), .B(n3886), .Z(n1918) );
  AN2 U1748 ( .A(n3882), .B(n495), .Z(n3886) );
  AN2 U1749 ( .A(n433), .B(n3883), .Z(n3882) );
  AN2 U1750 ( .A(ENCODER_CONTROL_IN[1]), .B(n385), .Z(n3883) );
  IV U1751 ( .A(n2591), .Z(U3_n725) );
  OR2 U1752 ( .A(n2593), .B(n3887), .Z(n2591) );
  OR2 U1753 ( .A(n1766), .B(n1765), .Z(n3887) );
  OR2 U1754 ( .A(n2595), .B(n3888), .Z(n2593) );
  OR2 U1755 ( .A(n1768), .B(n1767), .Z(n3888) );
  OR2 U1756 ( .A(n2597), .B(n3889), .Z(n2595) );
  OR2 U1757 ( .A(n1770), .B(n1769), .Z(n3889) );
  OR2 U1758 ( .A(n1771), .B(n3890), .Z(n2597) );
  OR2 U1759 ( .A(n1944), .B(n1772), .Z(n3890) );
  OR2 U1760 ( .A(n3891), .B(n3892), .Z(U29_Z_1) );
  OR2 U1761 ( .A(n3893), .B(n3894), .Z(n3892) );
  AN2 U1762 ( .A(n305), .B(ENCODER_DATA_IN[15]), .Z(n3894) );
  AN2 U1763 ( .A(ENCODER_DATA_IN[23]), .B(U34_CONTROL2), .Z(n3893) );
  OR2 U1764 ( .A(U33_CONTROL5), .B(n3895), .Z(n3891) );
  AN2 U1765 ( .A(U29_DATA1_1), .B(U29_CONTROL1), .Z(n3895) );
  OR2 U1766 ( .A(n3896), .B(n3897), .Z(U29_Z_0) );
  OR2 U1767 ( .A(n3898), .B(n3899), .Z(n3897) );
  AN2 U1768 ( .A(ENCODER_DATA_IN[22]), .B(U34_CONTROL2), .Z(n3899) );
  AN2 U1769 ( .A(U29_DATA1_0), .B(U29_CONTROL1), .Z(n3898) );
  AN2 U1770 ( .A(n305), .B(ENCODER_DATA_IN[14]), .Z(n3896) );
  OR2 U1771 ( .A(n3900), .B(n3901), .Z(U29_DATA1_1) );
  OR2 U1772 ( .A(n1905), .B(n1902), .Z(n3900) );
  OR2 U1773 ( .A(n3902), .B(n3903), .Z(U29_DATA1_0) );
  OR2 U1774 ( .A(n3904), .B(n3905), .Z(U28_Z_2) );
  OR2 U1775 ( .A(n3906), .B(n3907), .Z(n3905) );
  AN2 U1776 ( .A(ENCODER_DATA_IN[26]), .B(U34_CONTROL2), .Z(n3907) );
  AN2 U1777 ( .A(ENCODER_DATA_IN[18]), .B(U28_CONTROL4), .Z(n3906) );
  OR2 U1778 ( .A(U33_CONTROL5), .B(n3908), .Z(n3904) );
  AN2 U1779 ( .A(U28_DATA1_2), .B(U29_CONTROL1), .Z(n3908) );
  OR2 U1780 ( .A(n3909), .B(n3910), .Z(U28_Z_1) );
  OR2 U1781 ( .A(n3911), .B(n3912), .Z(n3910) );
  AN2 U1782 ( .A(ENCODER_DATA_IN[25]), .B(U34_CONTROL2), .Z(n3912) );
  AN2 U1783 ( .A(ENCODER_DATA_IN[17]), .B(U28_CONTROL4), .Z(n3911) );
  OR2 U1784 ( .A(U33_CONTROL5), .B(n3913), .Z(n3909) );
  AN2 U1785 ( .A(U28_DATA1_1), .B(U29_CONTROL1), .Z(n3913) );
  OR2 U1786 ( .A(n3914), .B(n3915), .Z(U28_Z_0) );
  OR2 U1787 ( .A(n3916), .B(n3917), .Z(n3915) );
  AN2 U1788 ( .A(ENCODER_DATA_IN[24]), .B(U34_CONTROL2), .Z(n3917) );
  AN2 U1789 ( .A(ENCODER_DATA_IN[16]), .B(U28_CONTROL4), .Z(n3916) );
  OR2 U1790 ( .A(U33_CONTROL5), .B(n3918), .Z(n3914) );
  AN2 U1791 ( .A(U28_DATA1_0), .B(U29_CONTROL1), .Z(n3918) );
  OR2 U1792 ( .A(n3919), .B(n3920), .Z(U28_DATA1_2) );
  OR2 U1793 ( .A(n1904), .B(n1902), .Z(n3919) );
  OR2 U1794 ( .A(n3921), .B(n3920), .Z(U28_DATA1_1) );
  OR2 U1795 ( .A(n1900), .B(n3922), .Z(n3920) );
  OR2 U1796 ( .A(n1905), .B(n1903), .Z(n3921) );
  OR2 U1797 ( .A(n3923), .B(n3901), .Z(U28_DATA1_0) );
  OR2 U1798 ( .A(n1901), .B(n3922), .Z(n3901) );
  OR2 U1799 ( .A(n1899), .B(n1913), .Z(n3922) );
  IV U1800 ( .A(n3924), .Z(n1913) );
  OR2 U1801 ( .A(n3925), .B(n3926), .Z(n3924) );
  OR2 U1802 ( .A(n3927), .B(n3928), .Z(n3926) );
  OR2 U1803 ( .A(n391), .B(n390), .Z(n3928) );
  OR2 U1804 ( .A(n510), .B(n447), .Z(n3927) );
  OR2 U1805 ( .A(n3929), .B(n3930), .Z(n3925) );
  OR2 U1806 ( .A(n630), .B(n572), .Z(n3930) );
  OR2 U1807 ( .A(n692), .B(n3931), .Z(n3929) );
  OR2 U1808 ( .A(n808), .B(n746), .Z(n3931) );
  AN2 U1809 ( .A(n808), .B(n3932), .Z(n1899) );
  AN2 U1810 ( .A(n3933), .B(n747), .Z(n3932) );
  OR2 U1811 ( .A(n1904), .B(n1903), .Z(n3923) );
  OR2 U1812 ( .A(n3934), .B(n3935), .Z(U27_Z_1) );
  OR2 U1813 ( .A(n3936), .B(n3937), .Z(n3935) );
  AN2 U1814 ( .A(ENCODER_DATA_IN[20]), .B(U28_CONTROL4), .Z(n3937) );
  AN2 U1815 ( .A(U27_DATA1_1), .B(U29_CONTROL1), .Z(n3936) );
  AN2 U1816 ( .A(ENCODER_DATA_IN[28]), .B(U34_CONTROL2), .Z(n3934) );
  OR2 U1817 ( .A(n3938), .B(n3939), .Z(U27_Z_0) );
  OR2 U1818 ( .A(n3940), .B(n3941), .Z(n3939) );
  AN2 U1819 ( .A(ENCODER_DATA_IN[19]), .B(U28_CONTROL4), .Z(n3941) );
  AN2 U1820 ( .A(U27_DATA1_0), .B(U29_CONTROL1), .Z(n3940) );
  OR2 U1821 ( .A(n1535), .B(U32_CONTROL1), .Z(U29_CONTROL1) );
  OR2 U1822 ( .A(n1551), .B(U34_CONTROL1), .Z(U32_CONTROL1) );
  OR2 U1823 ( .A(n1663), .B(n2579), .Z(U34_CONTROL1) );
  AN2 U1824 ( .A(ENCODER_DATA_IN[27]), .B(U34_CONTROL2), .Z(n3938) );
  OR2 U1825 ( .A(n3902), .B(n3942), .Z(U27_DATA1_1) );
  OR2 U1826 ( .A(n1905), .B(n1904), .Z(n3902) );
  AN2 U1827 ( .A(n3943), .B(n510), .Z(n1904) );
  AN2 U1828 ( .A(n447), .B(n3944), .Z(n1905) );
  OR2 U1829 ( .A(n3903), .B(n3942), .Z(U27_DATA1_0) );
  OR2 U1830 ( .A(n1901), .B(n1900), .Z(n3942) );
  AN2 U1831 ( .A(n3933), .B(n746), .Z(n1900) );
  AN2 U1832 ( .A(n3945), .B(n693), .Z(n3933) );
  AN2 U1833 ( .A(n692), .B(n3945), .Z(n1901) );
  AN2 U1834 ( .A(n631), .B(n3946), .Z(n3945) );
  OR2 U1835 ( .A(n1903), .B(n1902), .Z(n3903) );
  AN2 U1836 ( .A(n3946), .B(n630), .Z(n1902) );
  AN2 U1837 ( .A(n573), .B(n3947), .Z(n3946) );
  AN2 U1838 ( .A(n572), .B(n3947), .Z(n1903) );
  AN2 U1839 ( .A(n3943), .B(n511), .Z(n3947) );
  AN2 U1840 ( .A(n448), .B(n3944), .Z(n3943) );
  AN2 U1841 ( .A(ENCODER_CONTROL_IN[2]), .B(n392), .Z(n3944) );
  OR2 U1842 ( .A(n3948), .B(n3949), .Z(U26_Z_2) );
  OR2 U1843 ( .A(n3950), .B(n3951), .Z(n3949) );
  AN2 U1844 ( .A(ENCODER_DATA_IN[31]), .B(U34_CONTROL2), .Z(n3951) );
  AN2 U1845 ( .A(ENCODER_DATA_IN[23]), .B(U28_CONTROL4), .Z(n3950) );
  OR2 U1846 ( .A(U33_CONTROL5), .B(n3952), .Z(n3948) );
  AN2 U1847 ( .A(n301), .B(U26_DATA1_2), .Z(n3952) );
  OR2 U1848 ( .A(n3953), .B(n3954), .Z(U26_Z_1) );
  OR2 U1849 ( .A(n3955), .B(n3956), .Z(n3954) );
  AN2 U1850 ( .A(ENCODER_DATA_IN[30]), .B(U34_CONTROL2), .Z(n3956) );
  AN2 U1851 ( .A(ENCODER_DATA_IN[22]), .B(U28_CONTROL4), .Z(n3955) );
  OR2 U1852 ( .A(U33_CONTROL5), .B(n3957), .Z(n3953) );
  AN2 U1853 ( .A(n301), .B(U26_DATA1_1), .Z(n3957) );
  OR2 U1854 ( .A(n3958), .B(n3959), .Z(U26_Z_0) );
  OR2 U1855 ( .A(n3960), .B(n3961), .Z(n3959) );
  AN2 U1856 ( .A(ENCODER_DATA_IN[21]), .B(U28_CONTROL4), .Z(n3961) );
  OR2 U1857 ( .A(n1503), .B(U25_CONTROL5), .Z(U28_CONTROL4) );
  AN2 U1858 ( .A(n301), .B(U26_DATA1_0), .Z(n3960) );
  AN2 U1859 ( .A(ENCODER_DATA_IN[29]), .B(U34_CONTROL2), .Z(n3958) );
  OR2 U1860 ( .A(n1583), .B(U25_CONTROL2), .Z(U34_CONTROL2) );
  OR2 U1861 ( .A(n3962), .B(n3963), .Z(U26_DATA1_2) );
  OR2 U1862 ( .A(n1889), .B(n1888), .Z(n3962) );
  OR2 U1863 ( .A(n3964), .B(n3963), .Z(U26_DATA1_1) );
  OR2 U1864 ( .A(n1886), .B(n3965), .Z(n3963) );
  OR2 U1865 ( .A(n1890), .B(n1887), .Z(n3964) );
  OR2 U1866 ( .A(n3966), .B(n3967), .Z(U26_DATA1_0) );
  OR2 U1867 ( .A(n3968), .B(n3969), .Z(U25_Z_1) );
  OR2 U1868 ( .A(n3970), .B(n3971), .Z(n3969) );
  AN2 U1869 ( .A(n1583), .B(ENCODER_DATA_IN[33]), .Z(n3971) );
  AN2 U1870 ( .A(ENCODER_DATA_IN[25]), .B(U25_CONTROL5), .Z(n3970) );
  OR2 U1871 ( .A(n3972), .B(n3973), .Z(n3968) );
  AN2 U1872 ( .A(n301), .B(U25_DATA1_1), .Z(n3972) );
  OR2 U1873 ( .A(n3974), .B(n3975), .Z(U25_Z_0) );
  OR2 U1874 ( .A(n3976), .B(n3977), .Z(n3975) );
  AN2 U1875 ( .A(n1583), .B(ENCODER_DATA_IN[32]), .Z(n3977) );
  AN2 U1876 ( .A(ENCODER_DATA_IN[24]), .B(U25_CONTROL5), .Z(n3976) );
  OR2 U1877 ( .A(n3978), .B(n3973), .Z(n3974) );
  OR2 U1878 ( .A(U33_CONTROL5), .B(n3979), .Z(n3973) );
  AN2 U1879 ( .A(n301), .B(U25_DATA1_0), .Z(n3978) );
  OR2 U1880 ( .A(n3980), .B(n3981), .Z(U25_DATA1_1) );
  OR2 U1881 ( .A(n1889), .B(n1887), .Z(n3980) );
  OR2 U1882 ( .A(n3982), .B(n3981), .Z(U25_DATA1_0) );
  OR2 U1883 ( .A(n1885), .B(n3965), .Z(n3981) );
  OR2 U1884 ( .A(n1884), .B(n1898), .Z(n3965) );
  IV U1885 ( .A(n3983), .Z(n1898) );
  OR2 U1886 ( .A(n3984), .B(n3985), .Z(n3983) );
  OR2 U1887 ( .A(n3986), .B(n3987), .Z(n3985) );
  OR2 U1888 ( .A(n398), .B(n397), .Z(n3987) );
  OR2 U1889 ( .A(n518), .B(n455), .Z(n3986) );
  OR2 U1890 ( .A(n3988), .B(n3989), .Z(n3984) );
  OR2 U1891 ( .A(n638), .B(n579), .Z(n3989) );
  OR2 U1892 ( .A(n699), .B(n3990), .Z(n3988) );
  OR2 U1893 ( .A(n823), .B(n752), .Z(n3990) );
  AN2 U1894 ( .A(n823), .B(n3991), .Z(n1884) );
  AN2 U1895 ( .A(n3992), .B(n753), .Z(n3991) );
  OR2 U1896 ( .A(n1890), .B(n1888), .Z(n3982) );
  OR2 U1897 ( .A(n3993), .B(n3994), .Z(U24_Z_1) );
  OR2 U1898 ( .A(n3995), .B(n3996), .Z(n3994) );
  AN2 U1899 ( .A(n1583), .B(ENCODER_DATA_IN[35]), .Z(n3996) );
  AN2 U1900 ( .A(ENCODER_DATA_IN[27]), .B(U25_CONTROL5), .Z(n3995) );
  OR2 U1901 ( .A(n3979), .B(n3997), .Z(n3993) );
  AN2 U1902 ( .A(n301), .B(U24_DATA1_1), .Z(n3997) );
  OR2 U1903 ( .A(n3998), .B(n3999), .Z(U24_Z_0) );
  OR2 U1904 ( .A(n4000), .B(n4001), .Z(n3999) );
  AN2 U1905 ( .A(n1583), .B(ENCODER_DATA_IN[34]), .Z(n4001) );
  AN2 U1906 ( .A(ENCODER_DATA_IN[26]), .B(U25_CONTROL5), .Z(n4000) );
  OR2 U1907 ( .A(n3979), .B(n4002), .Z(n3998) );
  AN2 U1908 ( .A(n301), .B(U24_DATA1_0), .Z(n4002) );
  AN2 U1909 ( .A(U25_CONTROL2), .B(n1805), .Z(n3979) );
  OR2 U1910 ( .A(n1567), .B(n2568), .Z(U25_CONTROL2) );
  OR2 U1911 ( .A(n3966), .B(n4003), .Z(U24_DATA1_1) );
  OR2 U1912 ( .A(n1890), .B(n1889), .Z(n3966) );
  AN2 U1913 ( .A(n4004), .B(n518), .Z(n1889) );
  AN2 U1914 ( .A(n455), .B(n4005), .Z(n1890) );
  OR2 U1915 ( .A(n3967), .B(n4003), .Z(U24_DATA1_0) );
  OR2 U1916 ( .A(n1886), .B(n1885), .Z(n4003) );
  AN2 U1917 ( .A(n3992), .B(n752), .Z(n1885) );
  AN2 U1918 ( .A(n4006), .B(n700), .Z(n3992) );
  AN2 U1919 ( .A(n699), .B(n4006), .Z(n1886) );
  AN2 U1920 ( .A(n639), .B(n4007), .Z(n4006) );
  OR2 U1921 ( .A(n1888), .B(n1887), .Z(n3967) );
  AN2 U1922 ( .A(n4007), .B(n638), .Z(n1887) );
  AN2 U1923 ( .A(n580), .B(n4008), .Z(n4007) );
  AN2 U1924 ( .A(n579), .B(n4008), .Z(n1888) );
  AN2 U1925 ( .A(n4004), .B(n519), .Z(n4008) );
  AN2 U1926 ( .A(n456), .B(n4005), .Z(n4004) );
  AN2 U1927 ( .A(ENCODER_CONTROL_IN[3]), .B(n399), .Z(n4005) );
  OR2 U1928 ( .A(n4009), .B(n4010), .Z(U23_Z_0) );
  OR2 U1929 ( .A(n4011), .B(n4012), .Z(n4010) );
  AN2 U1930 ( .A(n1583), .B(ENCODER_DATA_IN[36]), .Z(n4011) );
  OR2 U1931 ( .A(n4013), .B(n4014), .Z(n4009) );
  AN2 U1932 ( .A(ENCODER_DATA_IN[28]), .B(U25_CONTROL5), .Z(n4014) );
  AN2 U1933 ( .A(n296), .B(U23_DATA1_0), .Z(n4013) );
  OR2 U1934 ( .A(n4015), .B(n4016), .Z(U23_DATA1_0) );
  OR2 U1937 ( .A(n4018), .B(n4019), .Z(U20_Z_2) );
  OR2 U1938 ( .A(n4020), .B(n4021), .Z(n4019) );
  AN2 U1939 ( .A(n1583), .B(ENCODER_DATA_IN[39]), .Z(n4020) );
  OR2 U1940 ( .A(n4022), .B(n4023), .Z(n4018) );
  AN2 U1941 ( .A(ENCODER_DATA_IN[31]), .B(U25_CONTROL5), .Z(n4023) );
  AN2 U1942 ( .A(n296), .B(U20_DATA1_2), .Z(n4022) );
  OR2 U1943 ( .A(n4024), .B(n4025), .Z(U20_Z_1) );
  OR2 U1944 ( .A(n4026), .B(n4021), .Z(n4025) );
  AN2 U1945 ( .A(n1583), .B(ENCODER_DATA_IN[38]), .Z(n4026) );
  OR2 U1946 ( .A(n4027), .B(n4028), .Z(n4024) );
  AN2 U1947 ( .A(ENCODER_DATA_IN[30]), .B(U25_CONTROL5), .Z(n4028) );
  AN2 U1948 ( .A(n296), .B(U20_DATA1_1), .Z(n4027) );
  OR2 U1949 ( .A(n4029), .B(n4030), .Z(U20_Z_0) );
  OR2 U1950 ( .A(n4031), .B(n4021), .Z(n4030) );
  OR2 U1951 ( .A(n4012), .B(U33_CONTROL5), .Z(n4021) );
  AN2 U1952 ( .A(n295), .B(n1801), .Z(n4012) );
  AN2 U1953 ( .A(n1583), .B(ENCODER_DATA_IN[37]), .Z(n4031) );
  OR2 U1954 ( .A(n4032), .B(n4033), .Z(n4029) );
  AN2 U1955 ( .A(ENCODER_DATA_IN[29]), .B(U25_CONTROL5), .Z(n4033) );
  OR2 U1956 ( .A(n1487), .B(U19_CONTROL4), .Z(U25_CONTROL5) );
  AN2 U1957 ( .A(n296), .B(U20_DATA1_0), .Z(n4032) );
  OR2 U1958 ( .A(n4034), .B(n4035), .Z(U20_DATA1_2) );
  OR2 U1959 ( .A(n1875), .B(n1873), .Z(n4034) );
  OR2 U1960 ( .A(n4036), .B(n4037), .Z(U20_DATA1_1) );
  OR2 U1961 ( .A(n1874), .B(n1873), .Z(n4036) );
  OR2 U1962 ( .A(n4038), .B(n4037), .Z(U20_DATA1_0) );
  OR2 U1963 ( .A(n1871), .B(n4039), .Z(n4037) );
  OR2 U1964 ( .A(n1875), .B(n1872), .Z(n4038) );
  OR2 U1965 ( .A(n4040), .B(n4041), .Z(U19_Z_0) );
  OR2 U1966 ( .A(n4042), .B(n4043), .Z(n4041) );
  AN2 U1967 ( .A(ENCODER_DATA_IN[32]), .B(U19_CONTROL4), .Z(n4043) );
  AN2 U1968 ( .A(ENCODER_DATA_IN[40]), .B(U19_CONTROL2), .Z(n4042) );
  OR2 U1969 ( .A(U33_CONTROL5), .B(n4044), .Z(n4040) );
  AN2 U1970 ( .A(n296), .B(U19_DATA1_0), .Z(n4044) );
  OR2 U1971 ( .A(n4045), .B(n4035), .Z(U19_DATA1_0) );
  OR2 U1972 ( .A(n1870), .B(n4039), .Z(n4035) );
  OR2 U1973 ( .A(n1869), .B(n1883), .Z(n4039) );
  IV U1974 ( .A(n4046), .Z(n1883) );
  OR2 U1975 ( .A(n4047), .B(n4048), .Z(n4046) );
  OR2 U1976 ( .A(n4049), .B(n4050), .Z(n4048) );
  OR2 U1977 ( .A(n405), .B(n404), .Z(n4050) );
  OR2 U1978 ( .A(n526), .B(n463), .Z(n4049) );
  OR2 U1979 ( .A(n4051), .B(n4052), .Z(n4047) );
  OR2 U1980 ( .A(n646), .B(n586), .Z(n4052) );
  OR2 U1981 ( .A(n706), .B(n4053), .Z(n4051) );
  OR2 U1982 ( .A(n862), .B(n758), .Z(n4053) );
  AN2 U1983 ( .A(n862), .B(n4054), .Z(n1869) );
  AN2 U1984 ( .A(n4055), .B(n759), .Z(n4054) );
  OR2 U1985 ( .A(n1874), .B(n1872), .Z(n4045) );
  OR2 U1986 ( .A(n4056), .B(n4057), .Z(U18_Z_1) );
  OR2 U1987 ( .A(n4058), .B(n4059), .Z(n4057) );
  AN2 U1988 ( .A(ENCODER_DATA_IN[42]), .B(U19_CONTROL2), .Z(n4059) );
  AN2 U1989 ( .A(n296), .B(U18_DATA1_1), .Z(n4058) );
  AN2 U1990 ( .A(ENCODER_DATA_IN[34]), .B(U19_CONTROL4), .Z(n4056) );
  OR2 U1991 ( .A(n4060), .B(n4061), .Z(U18_Z_0) );
  OR2 U1992 ( .A(n4062), .B(n4063), .Z(n4061) );
  AN2 U1993 ( .A(ENCODER_DATA_IN[41]), .B(U19_CONTROL2), .Z(n4063) );
  AN2 U1994 ( .A(n296), .B(U18_DATA1_0), .Z(n4062) );
  AN2 U1995 ( .A(ENCODER_DATA_IN[33]), .B(U19_CONTROL4), .Z(n4060) );
  OR2 U1996 ( .A(n4015), .B(n4064), .Z(U18_DATA1_1) );
  OR2 U1997 ( .A(n1875), .B(n1874), .Z(n4015) );
  AN2 U1998 ( .A(n4065), .B(n526), .Z(n1874) );
  AN2 U1999 ( .A(n463), .B(n4066), .Z(n1875) );
  OR2 U2000 ( .A(n4016), .B(n4064), .Z(U18_DATA1_0) );
  OR2 U2001 ( .A(n1871), .B(n1870), .Z(n4064) );
  AN2 U2002 ( .A(n4055), .B(n758), .Z(n1870) );
  AN2 U2003 ( .A(n4067), .B(n707), .Z(n4055) );
  AN2 U2004 ( .A(n706), .B(n4067), .Z(n1871) );
  AN2 U2005 ( .A(n647), .B(n4068), .Z(n4067) );
  OR2 U2006 ( .A(n1873), .B(n1872), .Z(n4016) );
  AN2 U2007 ( .A(n4068), .B(n646), .Z(n1872) );
  AN2 U2008 ( .A(n587), .B(n4069), .Z(n4068) );
  AN2 U2009 ( .A(n586), .B(n4069), .Z(n1873) );
  AN2 U2010 ( .A(n4065), .B(n527), .Z(n4069) );
  AN2 U2011 ( .A(n464), .B(n4066), .Z(n4065) );
  AN2 U2012 ( .A(ENCODER_CONTROL_IN[4]), .B(n406), .Z(n4066) );
  OR2 U2013 ( .A(n4070), .B(n4071), .Z(U17_Z_4) );
  OR2 U2014 ( .A(n4072), .B(n4073), .Z(n4071) );
  AN2 U2015 ( .A(ENCODER_DATA_IN[39]), .B(U19_CONTROL4), .Z(n4073) );
  AN2 U2016 ( .A(ENCODER_DATA_IN[47]), .B(U19_CONTROL2), .Z(n4072) );
  OR2 U2017 ( .A(U33_CONTROL5), .B(n4074), .Z(n4070) );
  AN2 U2018 ( .A(n289), .B(U17_DATA1_4), .Z(n4074) );
  OR2 U2019 ( .A(n4075), .B(n4076), .Z(U17_Z_3) );
  OR2 U2020 ( .A(n4077), .B(n4078), .Z(n4076) );
  AN2 U2021 ( .A(ENCODER_DATA_IN[38]), .B(U19_CONTROL4), .Z(n4078) );
  AN2 U2022 ( .A(ENCODER_DATA_IN[46]), .B(U19_CONTROL2), .Z(n4077) );
  OR2 U2023 ( .A(U33_CONTROL5), .B(n4079), .Z(n4075) );
  AN2 U2024 ( .A(n289), .B(U17_DATA1_3), .Z(n4079) );
  OR2 U2025 ( .A(n4080), .B(n4081), .Z(U17_Z_2) );
  OR2 U2026 ( .A(n4082), .B(n4083), .Z(n4081) );
  AN2 U2027 ( .A(ENCODER_DATA_IN[37]), .B(U19_CONTROL4), .Z(n4083) );
  AN2 U2028 ( .A(ENCODER_DATA_IN[45]), .B(U19_CONTROL2), .Z(n4082) );
  OR2 U2029 ( .A(U33_CONTROL5), .B(n4084), .Z(n4080) );
  AN2 U2030 ( .A(n289), .B(U17_DATA1_2), .Z(n4084) );
  OR2 U2031 ( .A(n4085), .B(n4086), .Z(U17_Z_1) );
  OR2 U2032 ( .A(n4087), .B(n4088), .Z(n4086) );
  AN2 U2033 ( .A(ENCODER_DATA_IN[36]), .B(U19_CONTROL4), .Z(n4088) );
  AN2 U2034 ( .A(ENCODER_DATA_IN[44]), .B(U19_CONTROL2), .Z(n4087) );
  OR2 U2035 ( .A(U33_CONTROL5), .B(n4089), .Z(n4085) );
  AN2 U2036 ( .A(n289), .B(U17_DATA1_1), .Z(n4089) );
  OR2 U2037 ( .A(n4090), .B(n4091), .Z(U17_Z_0) );
  OR2 U2038 ( .A(n4092), .B(n4093), .Z(n4091) );
  AN2 U2039 ( .A(ENCODER_DATA_IN[43]), .B(U19_CONTROL2), .Z(n4093) );
  AN2 U2040 ( .A(n289), .B(U17_DATA1_0), .Z(n4092) );
  AN2 U2041 ( .A(ENCODER_DATA_IN[35]), .B(U19_CONTROL4), .Z(n4090) );
  OR2 U2042 ( .A(n1471), .B(n2560), .Z(U19_CONTROL4) );
  OR2 U2043 ( .A(n4094), .B(n4095), .Z(U17_DATA1_4) );
  OR2 U2044 ( .A(n1859), .B(n1857), .Z(n4094) );
  OR2 U2045 ( .A(n4096), .B(n4095), .Z(U17_DATA1_3) );
  OR2 U2046 ( .A(n1855), .B(n4097), .Z(n4095) );
  OR2 U2047 ( .A(n1860), .B(n1858), .Z(n4096) );
  OR2 U2048 ( .A(n4098), .B(n4099), .Z(U17_DATA1_2) );
  OR2 U2049 ( .A(n1859), .B(n1858), .Z(n4098) );
  OR2 U2050 ( .A(n4100), .B(n4099), .Z(U17_DATA1_1) );
  OR2 U2051 ( .A(n1856), .B(n4097), .Z(n4099) );
  OR2 U2052 ( .A(n1854), .B(n1868), .Z(n4097) );
  IV U2053 ( .A(n4101), .Z(n1868) );
  OR2 U2054 ( .A(n4102), .B(n4103), .Z(n4101) );
  OR2 U2055 ( .A(n4104), .B(n4105), .Z(n4103) );
  OR2 U2056 ( .A(n412), .B(n411), .Z(n4105) );
  OR2 U2057 ( .A(n534), .B(n470), .Z(n4104) );
  OR2 U2058 ( .A(n4106), .B(n4107), .Z(n4102) );
  OR2 U2059 ( .A(n654), .B(n593), .Z(n4107) );
  OR2 U2060 ( .A(n713), .B(n4108), .Z(n4106) );
  OR2 U2061 ( .A(n873), .B(n764), .Z(n4108) );
  AN2 U2062 ( .A(n873), .B(n4109), .Z(n1854) );
  AN2 U2063 ( .A(n4110), .B(n765), .Z(n4109) );
  OR2 U2064 ( .A(n1860), .B(n1857), .Z(n4100) );
  OR2 U2065 ( .A(n4111), .B(n4112), .Z(U17_DATA1_0) );
  OR2 U2066 ( .A(n4113), .B(n4114), .Z(U16_Z_1) );
  OR2 U2067 ( .A(n4115), .B(n4116), .Z(n4114) );
  AN2 U2068 ( .A(ENCODER_DATA_IN[49]), .B(U19_CONTROL2), .Z(n4116) );
  AN2 U2069 ( .A(n289), .B(U16_DATA1_1), .Z(n4115) );
  AN2 U2070 ( .A(ENCODER_DATA_IN[41]), .B(n309), .Z(n4113) );
  OR2 U2071 ( .A(n4117), .B(n4118), .Z(U16_Z_0) );
  OR2 U2072 ( .A(n4119), .B(n4120), .Z(n4118) );
  AN2 U2073 ( .A(ENCODER_DATA_IN[48]), .B(U19_CONTROL2), .Z(n4120) );
  AN2 U2074 ( .A(n289), .B(U16_DATA1_0), .Z(n4119) );
  AN2 U2075 ( .A(ENCODER_DATA_IN[40]), .B(n309), .Z(n4117) );
  OR2 U2076 ( .A(n4111), .B(n4121), .Z(U16_DATA1_1) );
  OR2 U2077 ( .A(n1860), .B(n1859), .Z(n4111) );
  AN2 U2078 ( .A(n4122), .B(n534), .Z(n1859) );
  AN2 U2079 ( .A(n470), .B(n4123), .Z(n1860) );
  OR2 U2080 ( .A(n4112), .B(n4121), .Z(U16_DATA1_0) );
  OR2 U2081 ( .A(n1856), .B(n1855), .Z(n4121) );
  AN2 U2082 ( .A(n4110), .B(n764), .Z(n1855) );
  AN2 U2083 ( .A(n4124), .B(n714), .Z(n4110) );
  AN2 U2084 ( .A(n713), .B(n4124), .Z(n1856) );
  AN2 U2085 ( .A(n655), .B(n4125), .Z(n4124) );
  OR2 U2086 ( .A(n1858), .B(n1857), .Z(n4112) );
  AN2 U2087 ( .A(n4125), .B(n654), .Z(n1857) );
  AN2 U2088 ( .A(n594), .B(n4126), .Z(n4125) );
  AN2 U2089 ( .A(n593), .B(n4126), .Z(n1858) );
  AN2 U2090 ( .A(n4122), .B(n535), .Z(n4126) );
  AN2 U2091 ( .A(n471), .B(n4123), .Z(n4122) );
  AN2 U2092 ( .A(ENCODER_CONTROL_IN[5]), .B(n413), .Z(n4123) );
  OR2 U2093 ( .A(n4127), .B(n4128), .Z(U15_Z_5) );
  OR2 U2094 ( .A(n4129), .B(n4130), .Z(n4128) );
  AN2 U2095 ( .A(ENCODER_DATA_IN[55]), .B(U19_CONTROL2), .Z(n4130) );
  AN2 U2096 ( .A(n286), .B(U15_DATA1_5), .Z(n4129) );
  AN2 U2097 ( .A(n309), .B(ENCODER_DATA_IN[47]), .Z(n4127) );
  OR2 U2098 ( .A(n4131), .B(n4132), .Z(U15_Z_4) );
  OR2 U2099 ( .A(n4133), .B(n4134), .Z(n4132) );
  AN2 U2100 ( .A(ENCODER_DATA_IN[46]), .B(n309), .Z(n4134) );
  AN2 U2101 ( .A(ENCODER_DATA_IN[54]), .B(U19_CONTROL2), .Z(n4133) );
  OR2 U2102 ( .A(U33_CONTROL5), .B(n4135), .Z(n4131) );
  AN2 U2103 ( .A(n286), .B(U15_DATA1_4), .Z(n4135) );
  OR2 U2104 ( .A(n4136), .B(n4137), .Z(U15_Z_3) );
  OR2 U2105 ( .A(n4138), .B(n4139), .Z(n4137) );
  AN2 U2106 ( .A(ENCODER_DATA_IN[45]), .B(n309), .Z(n4139) );
  AN2 U2107 ( .A(ENCODER_DATA_IN[53]), .B(U19_CONTROL2), .Z(n4138) );
  OR2 U2108 ( .A(U33_CONTROL5), .B(n4140), .Z(n4136) );
  AN2 U2109 ( .A(n286), .B(U15_DATA1_3), .Z(n4140) );
  OR2 U2110 ( .A(n4141), .B(n4142), .Z(U15_Z_2) );
  OR2 U2111 ( .A(n4143), .B(n4144), .Z(n4142) );
  AN2 U2112 ( .A(ENCODER_DATA_IN[44]), .B(n309), .Z(n4144) );
  AN2 U2113 ( .A(ENCODER_DATA_IN[52]), .B(U19_CONTROL2), .Z(n4143) );
  OR2 U2114 ( .A(U33_CONTROL5), .B(n4145), .Z(n4141) );
  AN2 U2115 ( .A(n286), .B(U15_DATA1_2), .Z(n4145) );
  OR2 U2116 ( .A(n4146), .B(n4147), .Z(U15_Z_1) );
  OR2 U2117 ( .A(n4148), .B(n4149), .Z(n4147) );
  AN2 U2118 ( .A(ENCODER_DATA_IN[43]), .B(n309), .Z(n4149) );
  AN2 U2119 ( .A(ENCODER_DATA_IN[51]), .B(U19_CONTROL2), .Z(n4148) );
  OR2 U2120 ( .A(U33_CONTROL5), .B(n4150), .Z(n4146) );
  AN2 U2121 ( .A(n286), .B(U15_DATA1_1), .Z(n4150) );
  OR2 U2122 ( .A(n4151), .B(n4152), .Z(U15_Z_0) );
  OR2 U2123 ( .A(n4153), .B(n4154), .Z(n4152) );
  AN2 U2124 ( .A(ENCODER_DATA_IN[50]), .B(U19_CONTROL2), .Z(n4154) );
  AN2 U2125 ( .A(n286), .B(U15_DATA1_0), .Z(n4153) );
  AN2 U2126 ( .A(ENCODER_DATA_IN[42]), .B(n309), .Z(n4151) );
  OR2 U2127 ( .A(n4155), .B(n4156), .Z(U15_DATA1_5) );
  OR2 U2128 ( .A(n4157), .B(n4158), .Z(U15_DATA1_4) );
  OR2 U2129 ( .A(n1844), .B(n1842), .Z(n4157) );
  OR2 U2130 ( .A(n4159), .B(n4158), .Z(U15_DATA1_3) );
  OR2 U2131 ( .A(n1840), .B(n4160), .Z(n4158) );
  OR2 U2132 ( .A(n1845), .B(n1843), .Z(n4159) );
  OR2 U2133 ( .A(n4161), .B(n4162), .Z(U15_DATA1_2) );
  OR2 U2134 ( .A(n1844), .B(n1843), .Z(n4161) );
  OR2 U2135 ( .A(n4163), .B(n4162), .Z(U15_DATA1_1) );
  OR2 U2136 ( .A(n1841), .B(n4160), .Z(n4162) );
  OR2 U2137 ( .A(n1839), .B(n1853), .Z(n4160) );
  IV U2138 ( .A(n4164), .Z(n1853) );
  OR2 U2139 ( .A(n4165), .B(n4166), .Z(n4164) );
  OR2 U2140 ( .A(n4167), .B(n4168), .Z(n4166) );
  OR2 U2141 ( .A(n426), .B(n425), .Z(n4168) );
  OR2 U2142 ( .A(n549), .B(n486), .Z(n4167) );
  OR2 U2143 ( .A(n4169), .B(n4170), .Z(n4165) );
  OR2 U2144 ( .A(n669), .B(n608), .Z(n4170) );
  OR2 U2145 ( .A(n726), .B(n4171), .Z(n4169) );
  OR2 U2146 ( .A(n888), .B(n781), .Z(n4171) );
  AN2 U2147 ( .A(n888), .B(n4172), .Z(n1839) );
  AN2 U2148 ( .A(n4173), .B(n782), .Z(n4172) );
  OR2 U2149 ( .A(n1845), .B(n1842), .Z(n4163) );
  OR2 U2150 ( .A(n4174), .B(n4155), .Z(U15_DATA1_0) );
  OR2 U2151 ( .A(n1843), .B(n1842), .Z(n4155) );
  AN2 U2152 ( .A(n4175), .B(n669), .Z(n1842) );
  AN2 U2153 ( .A(n608), .B(n4176), .Z(n1843) );
  OR2 U2154 ( .A(n4177), .B(n4178), .Z(U14_Z_0) );
  OR2 U2155 ( .A(n4179), .B(n4180), .Z(n4178) );
  AN2 U2156 ( .A(ENCODER_DATA_IN[56]), .B(U19_CONTROL2), .Z(n4180) );
  AN2 U2157 ( .A(n286), .B(U14_DATA1_0), .Z(n4179) );
  AN2 U2158 ( .A(ENCODER_DATA_IN[48]), .B(n1439), .Z(n4177) );
  OR2 U2159 ( .A(n4174), .B(n4156), .Z(U14_DATA1_0) );
  OR2 U2160 ( .A(n1841), .B(n1840), .Z(n4156) );
  AN2 U2161 ( .A(n4173), .B(n781), .Z(n1840) );
  AN2 U2162 ( .A(n4181), .B(n727), .Z(n4173) );
  AN2 U2163 ( .A(n726), .B(n4181), .Z(n1841) );
  AN2 U2164 ( .A(n670), .B(n4175), .Z(n4181) );
  AN2 U2165 ( .A(n609), .B(n4176), .Z(n4175) );
  AN2 U2166 ( .A(n4182), .B(n550), .Z(n4176) );
  OR2 U2167 ( .A(n1845), .B(n1844), .Z(n4174) );
  AN2 U2168 ( .A(n4182), .B(n549), .Z(n1844) );
  AN2 U2169 ( .A(n487), .B(n4183), .Z(n4182) );
  AN2 U2170 ( .A(n486), .B(n4183), .Z(n1845) );
  AN2 U2171 ( .A(ENCODER_CONTROL_IN[6]), .B(n427), .Z(n4183) );
  OR2 U2172 ( .A(n4184), .B(n4185), .Z(U13_Z_6) );
  OR2 U2173 ( .A(n4186), .B(n4187), .Z(n4185) );
  AN2 U2174 ( .A(ENCODER_DATA_IN[63]), .B(U19_CONTROL2), .Z(n4187) );
  AN2 U2175 ( .A(n283), .B(U13_DATA1_6), .Z(n4186) );
  AN2 U2176 ( .A(n1439), .B(ENCODER_DATA_IN[55]), .Z(n4184) );
  OR2 U2177 ( .A(n4188), .B(n4189), .Z(U13_Z_5) );
  OR2 U2178 ( .A(n4190), .B(n4191), .Z(n4189) );
  AN2 U2179 ( .A(ENCODER_DATA_IN[62]), .B(U19_CONTROL2), .Z(n4191) );
  AN2 U2180 ( .A(n283), .B(U13_DATA1_5), .Z(n4190) );
  AN2 U2181 ( .A(ENCODER_DATA_IN[54]), .B(n1439), .Z(n4188) );
  OR2 U2182 ( .A(n4192), .B(n4193), .Z(U13_Z_4) );
  OR2 U2183 ( .A(n4194), .B(n4195), .Z(n4193) );
  AN2 U2184 ( .A(ENCODER_DATA_IN[53]), .B(n1439), .Z(n4195) );
  AN2 U2185 ( .A(ENCODER_DATA_IN[61]), .B(U19_CONTROL2), .Z(n4194) );
  OR2 U2186 ( .A(U33_CONTROL5), .B(n4196), .Z(n4192) );
  AN2 U2187 ( .A(n283), .B(U13_DATA1_4), .Z(n4196) );
  OR2 U2188 ( .A(n4197), .B(n4198), .Z(U13_Z_3) );
  OR2 U2189 ( .A(n4199), .B(n4200), .Z(n4198) );
  AN2 U2190 ( .A(ENCODER_DATA_IN[52]), .B(n1439), .Z(n4200) );
  AN2 U2191 ( .A(ENCODER_DATA_IN[60]), .B(U19_CONTROL2), .Z(n4199) );
  OR2 U2192 ( .A(U33_CONTROL5), .B(n4201), .Z(n4197) );
  AN2 U2193 ( .A(n283), .B(U13_DATA1_3), .Z(n4201) );
  OR2 U2194 ( .A(n4202), .B(n4203), .Z(U13_Z_2) );
  OR2 U2195 ( .A(n4204), .B(n4205), .Z(n4203) );
  AN2 U2196 ( .A(ENCODER_DATA_IN[51]), .B(n1439), .Z(n4205) );
  AN2 U2197 ( .A(ENCODER_DATA_IN[59]), .B(U19_CONTROL2), .Z(n4204) );
  OR2 U2198 ( .A(U33_CONTROL5), .B(n4206), .Z(n4202) );
  AN2 U2199 ( .A(n283), .B(U13_DATA1_2), .Z(n4206) );
  OR2 U2200 ( .A(n4207), .B(n4208), .Z(U13_Z_1) );
  OR2 U2201 ( .A(n4209), .B(n4210), .Z(n4208) );
  AN2 U2202 ( .A(ENCODER_DATA_IN[50]), .B(n1439), .Z(n4210) );
  AN2 U2203 ( .A(ENCODER_DATA_IN[58]), .B(U19_CONTROL2), .Z(n4209) );
  OR2 U2204 ( .A(U33_CONTROL5), .B(n4211), .Z(n4207) );
  AN2 U2205 ( .A(n283), .B(U13_DATA1_1), .Z(n4211) );
  IV U2206 ( .A(n4212), .Z(U33_CONTROL5) );
  OR2 U2207 ( .A(n4213), .B(n4214), .Z(n4212) );
  OR2 U2208 ( .A(n2560), .B(n4215), .Z(n4214) );
  OR2 U2209 ( .A(n329), .B(n310), .Z(n4215) );
  OR2 U2210 ( .A(n287), .B(n4216), .Z(n310) );
  OR2 U2211 ( .A(n1535), .B(n1519), .Z(n4216) );
  OR2 U2212 ( .A(n1471), .B(n2569), .Z(n287) );
  OR2 U2213 ( .A(n1487), .B(n1503), .Z(n2569) );
  OR2 U2214 ( .A(n2579), .B(n4217), .Z(n329) );
  OR2 U2215 ( .A(n1599), .B(n2563), .Z(n4217) );
  OR2 U2216 ( .A(n1551), .B(n1567), .Z(n2563) );
  OR2 U2217 ( .A(n1439), .B(n1455), .Z(n2560) );
  OR2 U2218 ( .A(n1583), .B(n4218), .Z(n4213) );
  OR2 U2219 ( .A(n1663), .B(n1615), .Z(n4218) );
  OR2 U2220 ( .A(n4219), .B(n4220), .Z(U13_Z_0) );
  OR2 U2221 ( .A(n4221), .B(n4222), .Z(n4220) );
  AN2 U2222 ( .A(ENCODER_DATA_IN[57]), .B(U19_CONTROL2), .Z(n4222) );
  OR2 U2223 ( .A(n2568), .B(n4223), .Z(U19_CONTROL2) );
  OR2 U2224 ( .A(n1583), .B(n2579), .Z(n4223) );
  OR2 U2225 ( .A(n1631), .B(n1647), .Z(n2579) );
  OR2 U2226 ( .A(n1599), .B(n1615), .Z(n2568) );
  AN2 U2227 ( .A(n283), .B(U13_DATA1_0), .Z(n4221) );
  AN2 U2228 ( .A(ENCODER_DATA_IN[49]), .B(n1439), .Z(n4219) );
  OR2 U2229 ( .A(n4224), .B(n4225), .Z(U13_DATA1_6) );
  OR2 U2230 ( .A(n4226), .B(n4225), .Z(U13_DATA1_5) );
  OR2 U2231 ( .A(n1826), .B(n1825), .Z(n4225) );
  OR2 U2232 ( .A(n4227), .B(n4228), .Z(U13_DATA1_4) );
  OR2 U2233 ( .A(n1829), .B(n1827), .Z(n4227) );
  OR2 U2234 ( .A(n4229), .B(n4228), .Z(U13_DATA1_3) );
  OR2 U2235 ( .A(n1825), .B(n4230), .Z(n4228) );
  AN2 U2236 ( .A(n4231), .B(n802), .Z(n1825) );
  OR2 U2237 ( .A(n1830), .B(n1828), .Z(n4229) );
  OR2 U2238 ( .A(n4232), .B(n4233), .Z(U13_DATA1_2) );
  OR2 U2239 ( .A(n1829), .B(n1828), .Z(n4232) );
  OR2 U2240 ( .A(n4234), .B(n4233), .Z(U13_DATA1_1) );
  OR2 U2241 ( .A(n1826), .B(n4230), .Z(n4233) );
  OR2 U2242 ( .A(n1824), .B(n1838), .Z(n4230) );
  IV U2243 ( .A(n4235), .Z(n1838) );
  OR2 U2244 ( .A(n4236), .B(n4237), .Z(n4235) );
  OR2 U2245 ( .A(n4238), .B(n4239), .Z(n4237) );
  OR2 U2246 ( .A(n441), .B(n440), .Z(n4239) );
  OR2 U2247 ( .A(n564), .B(n502), .Z(n4238) );
  OR2 U2248 ( .A(n4240), .B(n4241), .Z(n4236) );
  OR2 U2249 ( .A(n684), .B(n623), .Z(n4241) );
  OR2 U2250 ( .A(n739), .B(n4242), .Z(n4240) );
  OR2 U2251 ( .A(n903), .B(n802), .Z(n4242) );
  AN2 U2252 ( .A(n903), .B(n4243), .Z(n1824) );
  AN2 U2253 ( .A(n4231), .B(n803), .Z(n4243) );
  AN2 U2254 ( .A(n4244), .B(n740), .Z(n4231) );
  AN2 U2255 ( .A(n739), .B(n4244), .Z(n1826) );
  AN2 U2256 ( .A(n685), .B(n4245), .Z(n4244) );
  OR2 U2257 ( .A(n1830), .B(n1827), .Z(n4234) );
  OR2 U2258 ( .A(n4224), .B(n4226), .Z(U13_DATA1_0) );
  OR2 U2259 ( .A(n1828), .B(n1827), .Z(n4226) );
  AN2 U2260 ( .A(n4245), .B(n684), .Z(n1827) );
  AN2 U2261 ( .A(n624), .B(n4246), .Z(n4245) );
  AN2 U2262 ( .A(n623), .B(n4246), .Z(n1828) );
  AN2 U2263 ( .A(n4247), .B(n565), .Z(n4246) );
  OR2 U2264 ( .A(n1830), .B(n1829), .Z(n4224) );
  AN2 U2265 ( .A(n4247), .B(n564), .Z(n1829) );
  AN2 U2266 ( .A(n503), .B(n4248), .Z(n4247) );
  AN2 U2267 ( .A(n502), .B(n4248), .Z(n1830) );
  AN2 U2268 ( .A(ENCODER_CONTROL_IN[7]), .B(n442), .Z(n4248) );
  AN2 U2332 ( .A(n4304), .B(U4_DATA1_7), .Z(n1363) );
  AN2 U2333 ( .A(n4305), .B(n1971), .Z(n1297) );
  AN2 U2334 ( .A(n1970), .B(n4306), .Z(n4305) );
  IV U2335 ( .A(n1364), .Z(n4306) );
  AN2 U2336 ( .A(n4304), .B(n2460), .Z(n1296) );
  IV U2337 ( .A(n4307), .Z(n4304) );
  OR2 U2338 ( .A(n2491), .B(n4308), .Z(n4307) );
  OR2 U2339 ( .A(n1971), .B(n1364), .Z(n4308) );
  AN2 U2340 ( .A(n4309), .B(n4310), .Z(n1237) );
  AN2 U2341 ( .A(n4311), .B(n919), .Z(n4310) );
  AN2 U2342 ( .A(n1970), .B(n4312), .Z(n4311) );
  IV U2343 ( .A(n1046), .Z(n4312) );
  AN2 U2344 ( .A(n4313), .B(n949), .Z(n4309) );
  AN2 U2345 ( .A(n940), .B(n931), .Z(n4313) );
  AN2 U2346 ( .A(DATA_VALID), .B(n2491), .Z(n1062) );
  OR2 U2347 ( .A(n4314), .B(n4315), .Z(U6_Z_8) );
  AN2 U2348 ( .A(n4316), .B(n2412), .Z(n4315) );
  IV U2349 ( .A(U4_DATA1_8), .Z(n2412) );
  AN2 U2350 ( .A(n4317), .B(n4318), .Z(n4316) );
  AN2 U2351 ( .A(n4319), .B(U4_DATA1_7), .Z(n4317) );
  AN2 U2352 ( .A(n4320), .B(U4_DATA1_8), .Z(n4314) );
  OR2 U2353 ( .A(n4321), .B(n4322), .Z(n4320) );
  AN2 U2354 ( .A(n4318), .B(n2460), .Z(n4321) );
  OR2 U2355 ( .A(n4323), .B(n4324), .Z(U6_Z_7) );
  AN2 U2356 ( .A(n4325), .B(n2460), .Z(n4324) );
  IV U2357 ( .A(U4_DATA1_7), .Z(n2460) );
  AN2 U2358 ( .A(n4318), .B(n4319), .Z(n4325) );
  IV U2359 ( .A(n4326), .Z(n4319) );
  AN2 U2360 ( .A(n4322), .B(U4_DATA1_7), .Z(n4323) );
  OR2 U2361 ( .A(n4327), .B(n4328), .Z(n4322) );
  AN2 U2362 ( .A(n4318), .B(n4326), .Z(n4327) );
  OR2 U2363 ( .A(n4329), .B(n4330), .Z(n4326) );
  OR2 U2364 ( .A(n4331), .B(n4332), .Z(n4330) );
  OR2 U2365 ( .A(n4333), .B(n4334), .Z(U6_Z_6) );
  AN2 U2366 ( .A(n4335), .B(n4329), .Z(n4334) );
  IV U2367 ( .A(U4_DATA1_6), .Z(n4329) );
  AN2 U2368 ( .A(n4336), .B(n4318), .Z(n4335) );
  AN2 U2369 ( .A(U4_DATA1_5), .B(n4337), .Z(n4336) );
  AN2 U2370 ( .A(U4_DATA1_6), .B(n4338), .Z(n4333) );
  OR2 U2371 ( .A(n4339), .B(n4340), .Z(n4338) );
  AN2 U2372 ( .A(n4318), .B(n4332), .Z(n4339) );
  OR2 U2373 ( .A(n4341), .B(n4342), .Z(U6_Z_5) );
  AN2 U2374 ( .A(n4343), .B(n4332), .Z(n4342) );
  IV U2375 ( .A(U4_DATA1_5), .Z(n4332) );
  AN2 U2376 ( .A(n4318), .B(n4337), .Z(n4343) );
  IV U2377 ( .A(n4331), .Z(n4337) );
  AN2 U2378 ( .A(U4_DATA1_5), .B(n4340), .Z(n4341) );
  OR2 U2379 ( .A(n4344), .B(n4328), .Z(n4340) );
  AN2 U2380 ( .A(n4318), .B(n4331), .Z(n4344) );
  OR2 U2381 ( .A(n4345), .B(n4346), .Z(n4331) );
  OR2 U2382 ( .A(n4347), .B(n4348), .Z(n4346) );
  OR2 U2383 ( .A(n4349), .B(n4350), .Z(U6_Z_4) );
  AN2 U2384 ( .A(n4351), .B(n4345), .Z(n4350) );
  IV U2385 ( .A(U4_DATA1_4), .Z(n4345) );
  AN2 U2386 ( .A(n4352), .B(n4318), .Z(n4351) );
  AN2 U2387 ( .A(U4_DATA1_3), .B(n4353), .Z(n4352) );
  AN2 U2388 ( .A(U4_DATA1_4), .B(n4354), .Z(n4349) );
  OR2 U2389 ( .A(n4355), .B(n4356), .Z(n4354) );
  AN2 U2390 ( .A(n4318), .B(n4348), .Z(n4355) );
  OR2 U2391 ( .A(n4357), .B(n4358), .Z(U6_Z_3) );
  AN2 U2392 ( .A(n4359), .B(n4348), .Z(n4358) );
  IV U2393 ( .A(U4_DATA1_3), .Z(n4348) );
  AN2 U2394 ( .A(n4318), .B(n4353), .Z(n4359) );
  IV U2395 ( .A(n4347), .Z(n4353) );
  AN2 U2396 ( .A(U4_DATA1_3), .B(n4356), .Z(n4357) );
  OR2 U2397 ( .A(n4360), .B(n4328), .Z(n4356) );
  AN2 U2398 ( .A(n4318), .B(n4347), .Z(n4360) );
  OR2 U2399 ( .A(n4361), .B(n4362), .Z(n4347) );
  OR2 U2400 ( .A(n4363), .B(n4364), .Z(n4362) );
  OR2 U2401 ( .A(n4365), .B(n4366), .Z(U6_Z_2) );
  AN2 U2402 ( .A(n4367), .B(n4361), .Z(n4366) );
  IV U2403 ( .A(U4_DATA1_2), .Z(n4361) );
  AN2 U2404 ( .A(n4368), .B(n4318), .Z(n4367) );
  AN2 U2405 ( .A(U4_DATA1_1), .B(U4_DATA1_0), .Z(n4368) );
  AN2 U2406 ( .A(U4_DATA1_2), .B(n4369), .Z(n4365) );
  OR2 U2407 ( .A(n4370), .B(n4371), .Z(n4369) );
  AN2 U2408 ( .A(n4318), .B(n4364), .Z(n4370) );
  OR2 U2409 ( .A(n4372), .B(n4373), .Z(U6_Z_1) );
  AN2 U2410 ( .A(n4374), .B(n4364), .Z(n4373) );
  IV U2411 ( .A(U4_DATA1_1), .Z(n4364) );
  AN2 U2412 ( .A(n4318), .B(U4_DATA1_0), .Z(n4374) );
  AN2 U2413 ( .A(U4_DATA1_1), .B(n4371), .Z(n4372) );
  OR2 U2414 ( .A(n4375), .B(n4328), .Z(n4371) );
  OR2 U2415 ( .A(n4375), .B(n4376), .Z(U6_Z_0) );
  AN2 U2416 ( .A(n4328), .B(U4_DATA1_0), .Z(n4376) );
  AN2 U2417 ( .A(n4377), .B(n1046), .Z(n4328) );
  AN2 U2418 ( .A(n4318), .B(n4363), .Z(n4375) );
  IV U2419 ( .A(U4_DATA1_0), .Z(n4363) );
  AN2 U2420 ( .A(n4377), .B(DATA_VALID), .Z(n4318) );
  IV U2421 ( .A(n1057), .Z(n4377) );
  OR2 U2422 ( .A(n4378), .B(n4379), .Z(U5_Z_9) );
  OR2 U2423 ( .A(n4380), .B(n4381), .Z(n4379) );
  OR2 U2424 ( .A(n4382), .B(n4383), .Z(n4381) );
  AN2 U2425 ( .A(U7_DATA4_9), .B(n4384), .Z(n4383) );
  AN2 U2426 ( .A(U7_DATA6_9), .B(n4385), .Z(n4382) );
  AN2 U2427 ( .A(n2661), .B(U7_DATA1_9), .Z(n4380) );
  OR2 U2428 ( .A(n4386), .B(n4387), .Z(n4378) );
  OR2 U2429 ( .A(n4388), .B(n4389), .Z(n4387) );
  AN2 U2430 ( .A(n4390), .B(ENCODER_DATA_OUT[17]), .Z(n4389) );
  AN2 U2431 ( .A(TEST_PAT_SEED_A[9]), .B(n4391), .Z(n4388) );
  AN2 U2432 ( .A(TEST_PAT_SEED_B[9]), .B(n4392), .Z(n4386) );
  OR2 U2433 ( .A(n4393), .B(n4394), .Z(U5_Z_8) );
  OR2 U2434 ( .A(n4395), .B(n4396), .Z(n4394) );
  OR2 U2435 ( .A(n4397), .B(n4398), .Z(n4396) );
  AN2 U2436 ( .A(U7_DATA4_8), .B(n4384), .Z(n4398) );
  AN2 U2437 ( .A(U7_DATA6_8), .B(n4385), .Z(n4397) );
  AN2 U2438 ( .A(n2661), .B(U7_DATA1_8), .Z(n4395) );
  OR2 U2439 ( .A(n4399), .B(n4400), .Z(n4393) );
  OR2 U2440 ( .A(n4401), .B(n4402), .Z(n4400) );
  AN2 U2441 ( .A(n4390), .B(ENCODER_DATA_OUT[16]), .Z(n4402) );
  AN2 U2442 ( .A(TEST_PAT_SEED_A[8]), .B(n4391), .Z(n4401) );
  AN2 U2443 ( .A(TEST_PAT_SEED_B[8]), .B(n4392), .Z(n4399) );
  OR2 U2444 ( .A(n4403), .B(n4404), .Z(U5_Z_7) );
  OR2 U2445 ( .A(n4405), .B(n4406), .Z(n4404) );
  OR2 U2446 ( .A(n4407), .B(n4408), .Z(n4406) );
  AN2 U2447 ( .A(U7_DATA4_7), .B(n4384), .Z(n4408) );
  AN2 U2448 ( .A(U7_DATA6_7), .B(n4385), .Z(n4407) );
  AN2 U2449 ( .A(n2661), .B(U7_DATA1_7), .Z(n4405) );
  OR2 U2450 ( .A(n4409), .B(n4410), .Z(n4403) );
  OR2 U2451 ( .A(n4411), .B(n4412), .Z(n4410) );
  AN2 U2452 ( .A(n4390), .B(ENCODER_DATA_OUT[15]), .Z(n4412) );
  AN2 U2453 ( .A(TEST_PAT_SEED_A[7]), .B(n4391), .Z(n4411) );
  AN2 U2454 ( .A(TEST_PAT_SEED_B[7]), .B(n4392), .Z(n4409) );
  OR2 U2455 ( .A(n4413), .B(n4414), .Z(U5_Z_6) );
  OR2 U2456 ( .A(n4415), .B(n4416), .Z(n4414) );
  OR2 U2457 ( .A(n4417), .B(n4418), .Z(n4416) );
  AN2 U2458 ( .A(U7_DATA4_6), .B(n4384), .Z(n4418) );
  AN2 U2459 ( .A(U7_DATA6_6), .B(n4385), .Z(n4417) );
  AN2 U2460 ( .A(n2661), .B(U7_DATA1_6), .Z(n4415) );
  OR2 U2461 ( .A(n4419), .B(n4420), .Z(n4413) );
  OR2 U2462 ( .A(n4421), .B(n4422), .Z(n4420) );
  AN2 U2463 ( .A(n4390), .B(ENCODER_DATA_OUT[14]), .Z(n4422) );
  AN2 U2464 ( .A(TEST_PAT_SEED_A[6]), .B(n4391), .Z(n4421) );
  AN2 U2465 ( .A(TEST_PAT_SEED_B[6]), .B(n4392), .Z(n4419) );
  OR2 U2466 ( .A(n4423), .B(n4424), .Z(U5_Z_57) );
  OR2 U2467 ( .A(n4425), .B(n4426), .Z(n4424) );
  OR2 U2468 ( .A(n4427), .B(n4428), .Z(n4426) );
  AN2 U2469 ( .A(U7_DATA4_57), .B(n4384), .Z(n4428) );
  AN2 U2470 ( .A(U7_DATA6_57), .B(n4385), .Z(n4427) );
  AN2 U2471 ( .A(n2661), .B(U7_DATA1_57), .Z(n4425) );
  OR2 U2472 ( .A(n4429), .B(n4430), .Z(n4423) );
  OR2 U2473 ( .A(n4431), .B(n4432), .Z(n4430) );
  AN2 U2474 ( .A(ENCODER_DATA_OUT[65]), .B(n4390), .Z(n4432) );
  AN2 U2475 ( .A(n4433), .B(n4434), .Z(ENCODER_DATA_OUT[65]) );
  IV U2476 ( .A(n4435), .Z(n4434) );
  AN2 U2477 ( .A(n4436), .B(ENCODER_DATA_OUT[7]), .Z(n4435) );
  OR2 U2478 ( .A(ENCODER_DATA_OUT[7]), .B(n4436), .Z(n4433) );
  OR2 U2479 ( .A(n4437), .B(n4438), .Z(n4436) );
  AN2 U2480 ( .A(n4439), .B(n4440), .Z(n4438) );
  IV U2481 ( .A(n4441), .Z(n4437) );
  OR2 U2482 ( .A(n4440), .B(n4439), .Z(n4441) );
  OR2 U2483 ( .A(n4442), .B(n4443), .Z(n4440) );
  OR2 U2484 ( .A(n279), .B(n4444), .Z(n4443) );
  AN2 U2485 ( .A(ENCODER_DATA_IN[63]), .B(n4445), .Z(n4444) );
  AN2 U2486 ( .A(U13_Z_6), .B(n4446), .Z(n4442) );
  AN2 U2487 ( .A(TEST_PAT_SEED_A[57]), .B(n4391), .Z(n4431) );
  AN2 U2488 ( .A(TEST_PAT_SEED_B[57]), .B(n4392), .Z(n4429) );
  OR2 U2489 ( .A(n4447), .B(n4448), .Z(U5_Z_56) );
  OR2 U2490 ( .A(n4449), .B(n4450), .Z(n4448) );
  OR2 U2491 ( .A(n4451), .B(n4452), .Z(n4450) );
  AN2 U2492 ( .A(U7_DATA4_56), .B(n4384), .Z(n4452) );
  AN2 U2493 ( .A(U7_DATA6_56), .B(n4385), .Z(n4451) );
  AN2 U2494 ( .A(n2661), .B(U7_DATA1_56), .Z(n4449) );
  OR2 U2495 ( .A(n4453), .B(n4454), .Z(n4447) );
  OR2 U2496 ( .A(n4455), .B(n4456), .Z(n4454) );
  AN2 U2497 ( .A(ENCODER_DATA_OUT[64]), .B(n4390), .Z(n4456) );
  AN2 U2498 ( .A(n4457), .B(n4458), .Z(ENCODER_DATA_OUT[64]) );
  IV U2499 ( .A(n4459), .Z(n4458) );
  AN2 U2500 ( .A(n4460), .B(ENCODER_DATA_OUT[6]), .Z(n4459) );
  OR2 U2501 ( .A(ENCODER_DATA_OUT[6]), .B(n4460), .Z(n4457) );
  OR2 U2502 ( .A(n4461), .B(n4462), .Z(n4460) );
  IV U2503 ( .A(n4463), .Z(n4462) );
  OR2 U2504 ( .A(ENCODER_DATA_OUT[25]), .B(n4464), .Z(n4463) );
  AN2 U2505 ( .A(n4464), .B(ENCODER_DATA_OUT[25]), .Z(n4461) );
  IV U2506 ( .A(n4465), .Z(n4464) );
  OR2 U2507 ( .A(n4466), .B(n4467), .Z(n4465) );
  OR2 U2508 ( .A(n279), .B(n4468), .Z(n4467) );
  AN2 U2509 ( .A(ENCODER_DATA_IN[62]), .B(n4445), .Z(n4468) );
  AN2 U2510 ( .A(U13_Z_5), .B(n4446), .Z(n4466) );
  AN2 U2511 ( .A(TEST_PAT_SEED_A[56]), .B(n4391), .Z(n4455) );
  AN2 U2512 ( .A(TEST_PAT_SEED_B[56]), .B(n4392), .Z(n4453) );
  OR2 U2513 ( .A(n4469), .B(n4470), .Z(U5_Z_55) );
  OR2 U2514 ( .A(n4471), .B(n4472), .Z(n4470) );
  OR2 U2515 ( .A(n4473), .B(n4474), .Z(n4472) );
  AN2 U2516 ( .A(U7_DATA4_55), .B(n4384), .Z(n4474) );
  AN2 U2517 ( .A(U7_DATA6_55), .B(n4385), .Z(n4473) );
  AN2 U2518 ( .A(n2661), .B(U7_DATA1_55), .Z(n4471) );
  OR2 U2519 ( .A(n4475), .B(n4476), .Z(n4469) );
  OR2 U2520 ( .A(n4477), .B(n4478), .Z(n4476) );
  AN2 U2521 ( .A(ENCODER_DATA_OUT[63]), .B(n4390), .Z(n4478) );
  AN2 U2522 ( .A(n4479), .B(n4480), .Z(ENCODER_DATA_OUT[63]) );
  IV U2523 ( .A(n4481), .Z(n4480) );
  AN2 U2524 ( .A(n4482), .B(ENCODER_DATA_OUT[5]), .Z(n4481) );
  OR2 U2525 ( .A(ENCODER_DATA_OUT[5]), .B(n4482), .Z(n4479) );
  OR2 U2526 ( .A(n4483), .B(n4484), .Z(n4482) );
  IV U2527 ( .A(n4485), .Z(n4484) );
  OR2 U2528 ( .A(ENCODER_DATA_OUT[24]), .B(n4486), .Z(n4485) );
  AN2 U2529 ( .A(n4486), .B(ENCODER_DATA_OUT[24]), .Z(n4483) );
  IV U2530 ( .A(n4487), .Z(n4486) );
  OR2 U2531 ( .A(n4488), .B(n4489), .Z(n4487) );
  OR2 U2532 ( .A(n279), .B(n4490), .Z(n4489) );
  AN2 U2533 ( .A(ENCODER_DATA_IN[61]), .B(n4445), .Z(n4490) );
  AN2 U2534 ( .A(U13_Z_4), .B(n4446), .Z(n4488) );
  AN2 U2535 ( .A(TEST_PAT_SEED_A[55]), .B(n4391), .Z(n4477) );
  AN2 U2536 ( .A(TEST_PAT_SEED_B[55]), .B(n4392), .Z(n4475) );
  OR2 U2537 ( .A(n4491), .B(n4492), .Z(U5_Z_54) );
  OR2 U2538 ( .A(n4493), .B(n4494), .Z(n4492) );
  OR2 U2539 ( .A(n4495), .B(n4496), .Z(n4494) );
  AN2 U2540 ( .A(U7_DATA4_54), .B(n4384), .Z(n4496) );
  AN2 U2541 ( .A(U7_DATA6_54), .B(n4385), .Z(n4495) );
  AN2 U2542 ( .A(n2661), .B(U7_DATA1_54), .Z(n4493) );
  OR2 U2543 ( .A(n4497), .B(n4498), .Z(n4491) );
  OR2 U2544 ( .A(n4499), .B(n4500), .Z(n4498) );
  AN2 U2545 ( .A(ENCODER_DATA_OUT[62]), .B(n4390), .Z(n4500) );
  AN2 U2546 ( .A(n4501), .B(n4502), .Z(ENCODER_DATA_OUT[62]) );
  IV U2547 ( .A(n4503), .Z(n4502) );
  AN2 U2548 ( .A(n4504), .B(ENCODER_DATA_OUT[4]), .Z(n4503) );
  OR2 U2549 ( .A(ENCODER_DATA_OUT[4]), .B(n4504), .Z(n4501) );
  OR2 U2550 ( .A(n4505), .B(n4506), .Z(n4504) );
  IV U2551 ( .A(n4507), .Z(n4506) );
  OR2 U2552 ( .A(ENCODER_DATA_OUT[23]), .B(n4508), .Z(n4507) );
  AN2 U2553 ( .A(n4508), .B(ENCODER_DATA_OUT[23]), .Z(n4505) );
  IV U2554 ( .A(n4509), .Z(n4508) );
  OR2 U2555 ( .A(n4510), .B(n4511), .Z(n4509) );
  OR2 U2556 ( .A(n279), .B(n4512), .Z(n4511) );
  AN2 U2557 ( .A(ENCODER_DATA_IN[60]), .B(n4445), .Z(n4512) );
  AN2 U2558 ( .A(U13_Z_3), .B(n4446), .Z(n4510) );
  AN2 U2559 ( .A(TEST_PAT_SEED_A[54]), .B(n4391), .Z(n4499) );
  AN2 U2560 ( .A(TEST_PAT_SEED_B[54]), .B(n4392), .Z(n4497) );
  OR2 U2561 ( .A(n4513), .B(n4514), .Z(U5_Z_53) );
  OR2 U2562 ( .A(n4515), .B(n4516), .Z(n4514) );
  OR2 U2563 ( .A(n4517), .B(n4518), .Z(n4516) );
  AN2 U2564 ( .A(U7_DATA4_53), .B(n4384), .Z(n4518) );
  AN2 U2565 ( .A(U7_DATA6_53), .B(n4385), .Z(n4517) );
  AN2 U2566 ( .A(n2661), .B(U7_DATA1_53), .Z(n4515) );
  OR2 U2567 ( .A(n4519), .B(n4520), .Z(n4513) );
  OR2 U2568 ( .A(n4521), .B(n4522), .Z(n4520) );
  AN2 U2569 ( .A(ENCODER_DATA_OUT[61]), .B(n4390), .Z(n4522) );
  AN2 U2570 ( .A(n4523), .B(n4524), .Z(ENCODER_DATA_OUT[61]) );
  IV U2571 ( .A(n4525), .Z(n4524) );
  AN2 U2572 ( .A(n4526), .B(ENCODER_DATA_OUT[3]), .Z(n4525) );
  OR2 U2573 ( .A(ENCODER_DATA_OUT[3]), .B(n4526), .Z(n4523) );
  OR2 U2574 ( .A(n4527), .B(n4528), .Z(n4526) );
  IV U2575 ( .A(n4529), .Z(n4528) );
  OR2 U2576 ( .A(ENCODER_DATA_OUT[22]), .B(n4530), .Z(n4529) );
  AN2 U2577 ( .A(n4530), .B(ENCODER_DATA_OUT[22]), .Z(n4527) );
  IV U2578 ( .A(n4531), .Z(n4530) );
  OR2 U2579 ( .A(n4532), .B(n4533), .Z(n4531) );
  OR2 U2580 ( .A(n279), .B(n4534), .Z(n4533) );
  AN2 U2581 ( .A(ENCODER_DATA_IN[59]), .B(n4445), .Z(n4534) );
  AN2 U2582 ( .A(U13_Z_2), .B(n4446), .Z(n4532) );
  AN2 U2583 ( .A(TEST_PAT_SEED_A[53]), .B(n4391), .Z(n4521) );
  AN2 U2584 ( .A(TEST_PAT_SEED_B[53]), .B(n4392), .Z(n4519) );
  OR2 U2585 ( .A(n4535), .B(n4536), .Z(U5_Z_52) );
  OR2 U2586 ( .A(n4537), .B(n4538), .Z(n4536) );
  OR2 U2587 ( .A(n4539), .B(n4540), .Z(n4538) );
  AN2 U2588 ( .A(U7_DATA4_52), .B(n4384), .Z(n4540) );
  AN2 U2589 ( .A(U7_DATA6_52), .B(n4385), .Z(n4539) );
  AN2 U2590 ( .A(n2661), .B(U7_DATA1_52), .Z(n4537) );
  OR2 U2591 ( .A(n4541), .B(n4542), .Z(n4535) );
  OR2 U2592 ( .A(n4543), .B(n4544), .Z(n4542) );
  AN2 U2593 ( .A(ENCODER_DATA_OUT[60]), .B(n4390), .Z(n4544) );
  AN2 U2594 ( .A(n4545), .B(n4546), .Z(ENCODER_DATA_OUT[60]) );
  IV U2595 ( .A(n4547), .Z(n4546) );
  AN2 U2596 ( .A(n4548), .B(ENCODER_DATA_OUT[2]), .Z(n4547) );
  OR2 U2597 ( .A(ENCODER_DATA_OUT[2]), .B(n4548), .Z(n4545) );
  OR2 U2598 ( .A(n4549), .B(n4550), .Z(n4548) );
  IV U2599 ( .A(n4551), .Z(n4550) );
  OR2 U2600 ( .A(ENCODER_DATA_OUT[21]), .B(n4552), .Z(n4551) );
  AN2 U2601 ( .A(n4552), .B(ENCODER_DATA_OUT[21]), .Z(n4549) );
  IV U2602 ( .A(n4553), .Z(n4552) );
  OR2 U2603 ( .A(n4554), .B(n4555), .Z(n4553) );
  OR2 U2604 ( .A(n279), .B(n4556), .Z(n4555) );
  AN2 U2605 ( .A(ENCODER_DATA_IN[58]), .B(n4445), .Z(n4556) );
  AN2 U2606 ( .A(U13_Z_1), .B(n4446), .Z(n4554) );
  AN2 U2607 ( .A(TEST_PAT_SEED_A[52]), .B(n4391), .Z(n4543) );
  AN2 U2608 ( .A(TEST_PAT_SEED_B[52]), .B(n4392), .Z(n4541) );
  OR2 U2609 ( .A(n4557), .B(n4558), .Z(U5_Z_51) );
  OR2 U2610 ( .A(n4559), .B(n4560), .Z(n4558) );
  OR2 U2611 ( .A(n4561), .B(n4562), .Z(n4560) );
  AN2 U2612 ( .A(U7_DATA4_51), .B(n4384), .Z(n4562) );
  AN2 U2613 ( .A(U7_DATA6_51), .B(n4385), .Z(n4561) );
  AN2 U2614 ( .A(n2661), .B(U7_DATA1_51), .Z(n4559) );
  OR2 U2615 ( .A(n4563), .B(n4564), .Z(n4557) );
  OR2 U2616 ( .A(n4565), .B(n4566), .Z(n4564) );
  AN2 U2617 ( .A(n4390), .B(ENCODER_DATA_OUT[59]), .Z(n4566) );
  OR2 U2618 ( .A(n4567), .B(n4568), .Z(ENCODER_DATA_OUT[59]) );
  AN2 U2619 ( .A(n4569), .B(ENCODER_DATA_OUT[20]), .Z(n4568) );
  IV U2620 ( .A(n4570), .Z(n4567) );
  OR2 U2621 ( .A(ENCODER_DATA_OUT[20]), .B(n4569), .Z(n4570) );
  OR2 U2622 ( .A(n4571), .B(n4572), .Z(n4569) );
  AN2 U2623 ( .A(n4573), .B(n4574), .Z(n4572) );
  IV U2624 ( .A(n4575), .Z(n4573) );
  AN2 U2625 ( .A(U7_DATA1_57), .B(n4575), .Z(n4571) );
  OR2 U2626 ( .A(n4576), .B(n4577), .Z(n4575) );
  OR2 U2627 ( .A(n279), .B(n4578), .Z(n4577) );
  AN2 U2628 ( .A(ENCODER_DATA_IN[57]), .B(n4445), .Z(n4578) );
  AN2 U2629 ( .A(U13_Z_0), .B(n4446), .Z(n4576) );
  AN2 U2630 ( .A(TEST_PAT_SEED_A[51]), .B(n4391), .Z(n4565) );
  AN2 U2631 ( .A(TEST_PAT_SEED_B[51]), .B(n4392), .Z(n4563) );
  OR2 U2632 ( .A(n4579), .B(n4580), .Z(U5_Z_50) );
  OR2 U2633 ( .A(n4581), .B(n4582), .Z(n4580) );
  OR2 U2634 ( .A(n4583), .B(n4584), .Z(n4582) );
  AN2 U2635 ( .A(U7_DATA4_50), .B(n4384), .Z(n4584) );
  AN2 U2636 ( .A(U7_DATA6_50), .B(n4385), .Z(n4583) );
  AN2 U2637 ( .A(n2661), .B(U7_DATA1_50), .Z(n4581) );
  OR2 U2638 ( .A(n4585), .B(n4586), .Z(n4579) );
  OR2 U2639 ( .A(n4587), .B(n4588), .Z(n4586) );
  AN2 U2640 ( .A(n4390), .B(ENCODER_DATA_OUT[58]), .Z(n4588) );
  OR2 U2641 ( .A(n4589), .B(n4590), .Z(ENCODER_DATA_OUT[58]) );
  AN2 U2642 ( .A(n4591), .B(ENCODER_DATA_OUT[19]), .Z(n4590) );
  IV U2643 ( .A(n4592), .Z(n4589) );
  OR2 U2644 ( .A(ENCODER_DATA_OUT[19]), .B(n4591), .Z(n4592) );
  OR2 U2645 ( .A(n4593), .B(n4594), .Z(n4591) );
  AN2 U2646 ( .A(n4595), .B(n4596), .Z(n4594) );
  IV U2647 ( .A(n4597), .Z(n4595) );
  AN2 U2648 ( .A(U7_DATA1_56), .B(n4597), .Z(n4593) );
  OR2 U2649 ( .A(n4598), .B(n4599), .Z(n4597) );
  OR2 U2650 ( .A(n281), .B(n4600), .Z(n4599) );
  AN2 U2651 ( .A(ENCODER_DATA_IN[56]), .B(n4445), .Z(n4600) );
  AN2 U2652 ( .A(U14_Z_0), .B(n4446), .Z(n4598) );
  AN2 U2653 ( .A(TEST_PAT_SEED_A[50]), .B(n4391), .Z(n4587) );
  AN2 U2654 ( .A(TEST_PAT_SEED_B[50]), .B(n4392), .Z(n4585) );
  OR2 U2655 ( .A(n4601), .B(n4602), .Z(U5_Z_5) );
  OR2 U2656 ( .A(n4603), .B(n4604), .Z(n4602) );
  OR2 U2657 ( .A(n4605), .B(n4606), .Z(n4604) );
  AN2 U2658 ( .A(U7_DATA4_5), .B(n4384), .Z(n4606) );
  AN2 U2659 ( .A(U7_DATA6_5), .B(n4385), .Z(n4605) );
  AN2 U2660 ( .A(n2661), .B(U7_DATA1_5), .Z(n4603) );
  OR2 U2661 ( .A(n4607), .B(n4608), .Z(n4601) );
  OR2 U2662 ( .A(n4609), .B(n4610), .Z(n4608) );
  AN2 U2663 ( .A(n4390), .B(ENCODER_DATA_OUT[13]), .Z(n4610) );
  AN2 U2664 ( .A(TEST_PAT_SEED_A[5]), .B(n4391), .Z(n4609) );
  AN2 U2665 ( .A(TEST_PAT_SEED_B[5]), .B(n4392), .Z(n4607) );
  OR2 U2666 ( .A(n4611), .B(n4612), .Z(U5_Z_49) );
  OR2 U2667 ( .A(n4613), .B(n4614), .Z(n4612) );
  OR2 U2668 ( .A(n4615), .B(n4616), .Z(n4614) );
  AN2 U2669 ( .A(U7_DATA4_49), .B(n4384), .Z(n4616) );
  AN2 U2670 ( .A(U7_DATA6_49), .B(n4385), .Z(n4615) );
  AN2 U2671 ( .A(n2661), .B(U7_DATA1_49), .Z(n4613) );
  OR2 U2672 ( .A(n4617), .B(n4618), .Z(n4611) );
  OR2 U2673 ( .A(n4619), .B(n4620), .Z(n4618) );
  AN2 U2674 ( .A(n4390), .B(ENCODER_DATA_OUT[57]), .Z(n4620) );
  OR2 U2675 ( .A(n4621), .B(n4622), .Z(ENCODER_DATA_OUT[57]) );
  AN2 U2676 ( .A(n4623), .B(ENCODER_DATA_OUT[18]), .Z(n4622) );
  IV U2677 ( .A(n4624), .Z(n4621) );
  OR2 U2678 ( .A(ENCODER_DATA_OUT[18]), .B(n4623), .Z(n4624) );
  OR2 U2679 ( .A(n4625), .B(n4626), .Z(n4623) );
  AN2 U2680 ( .A(n4627), .B(n4628), .Z(n4626) );
  IV U2681 ( .A(n4629), .Z(n4627) );
  AN2 U2682 ( .A(U7_DATA1_55), .B(n4629), .Z(n4625) );
  OR2 U2683 ( .A(n4630), .B(n4631), .Z(n4629) );
  OR2 U2684 ( .A(n279), .B(n4632), .Z(n4631) );
  AN2 U2685 ( .A(ENCODER_DATA_IN[55]), .B(n4445), .Z(n4632) );
  AN2 U2686 ( .A(U15_Z_5), .B(n4446), .Z(n4630) );
  AN2 U2687 ( .A(TEST_PAT_SEED_A[49]), .B(n4391), .Z(n4619) );
  AN2 U2688 ( .A(TEST_PAT_SEED_B[49]), .B(n4392), .Z(n4617) );
  OR2 U2689 ( .A(n4633), .B(n4634), .Z(U5_Z_48) );
  OR2 U2690 ( .A(n4635), .B(n4636), .Z(n4634) );
  OR2 U2691 ( .A(n4637), .B(n4638), .Z(n4636) );
  AN2 U2692 ( .A(U7_DATA4_48), .B(n4384), .Z(n4638) );
  AN2 U2693 ( .A(U7_DATA6_48), .B(n4385), .Z(n4637) );
  AN2 U2694 ( .A(n2661), .B(U7_DATA1_48), .Z(n4635) );
  OR2 U2695 ( .A(n4639), .B(n4640), .Z(n4633) );
  OR2 U2696 ( .A(n4641), .B(n4642), .Z(n4640) );
  AN2 U2697 ( .A(n4390), .B(ENCODER_DATA_OUT[56]), .Z(n4642) );
  OR2 U2698 ( .A(n4643), .B(n4644), .Z(ENCODER_DATA_OUT[56]) );
  AN2 U2699 ( .A(n4645), .B(ENCODER_DATA_OUT[17]), .Z(n4644) );
  IV U2700 ( .A(n4646), .Z(n4643) );
  OR2 U2701 ( .A(ENCODER_DATA_OUT[17]), .B(n4645), .Z(n4646) );
  OR2 U2702 ( .A(n4647), .B(n4648), .Z(n4645) );
  AN2 U2703 ( .A(n4649), .B(n4650), .Z(n4648) );
  IV U2704 ( .A(n4651), .Z(n4649) );
  AN2 U2705 ( .A(U7_DATA1_54), .B(n4651), .Z(n4647) );
  OR2 U2706 ( .A(n4652), .B(n4653), .Z(n4651) );
  OR2 U2707 ( .A(n279), .B(n4654), .Z(n4653) );
  AN2 U2708 ( .A(ENCODER_DATA_IN[54]), .B(n4445), .Z(n4654) );
  AN2 U2709 ( .A(U15_Z_4), .B(n4446), .Z(n4652) );
  AN2 U2710 ( .A(n4655), .B(n4656), .Z(ENCODER_DATA_OUT[17]) );
  IV U2711 ( .A(n4657), .Z(n4656) );
  AN2 U2712 ( .A(n4658), .B(n4659), .Z(n4657) );
  OR2 U2713 ( .A(n4659), .B(n4658), .Z(n4655) );
  OR2 U2714 ( .A(n4660), .B(n4661), .Z(n4658) );
  AN2 U2715 ( .A(U7_DATA1_15), .B(n4662), .Z(n4661) );
  AN2 U2716 ( .A(U7_DATA1_34), .B(n4663), .Z(n4660) );
  IV U2717 ( .A(U7_DATA1_15), .Z(n4663) );
  OR2 U2718 ( .A(n4664), .B(n4665), .Z(n4659) );
  OR2 U2719 ( .A(n279), .B(n4666), .Z(n4665) );
  AN2 U2720 ( .A(ENCODER_DATA_IN[15]), .B(n4445), .Z(n4666) );
  AN2 U2721 ( .A(U32_Z_0), .B(n4446), .Z(n4664) );
  AN2 U2722 ( .A(TEST_PAT_SEED_A[48]), .B(n4391), .Z(n4641) );
  AN2 U2723 ( .A(TEST_PAT_SEED_B[48]), .B(n4392), .Z(n4639) );
  OR2 U2724 ( .A(n4667), .B(n4668), .Z(U5_Z_47) );
  OR2 U2725 ( .A(n4669), .B(n4670), .Z(n4668) );
  OR2 U2726 ( .A(n4671), .B(n4672), .Z(n4670) );
  AN2 U2727 ( .A(U7_DATA4_47), .B(n4384), .Z(n4672) );
  AN2 U2728 ( .A(U7_DATA6_47), .B(n4385), .Z(n4671) );
  AN2 U2729 ( .A(n2661), .B(U7_DATA1_47), .Z(n4669) );
  OR2 U2730 ( .A(n4673), .B(n4674), .Z(n4667) );
  OR2 U2731 ( .A(n4675), .B(n4676), .Z(n4674) );
  AN2 U2732 ( .A(n4390), .B(ENCODER_DATA_OUT[55]), .Z(n4676) );
  OR2 U2733 ( .A(n4677), .B(n4678), .Z(ENCODER_DATA_OUT[55]) );
  AN2 U2734 ( .A(n4679), .B(ENCODER_DATA_OUT[16]), .Z(n4678) );
  IV U2735 ( .A(n4680), .Z(n4677) );
  OR2 U2736 ( .A(ENCODER_DATA_OUT[16]), .B(n4679), .Z(n4680) );
  OR2 U2737 ( .A(n4681), .B(n4682), .Z(n4679) );
  AN2 U2738 ( .A(n4683), .B(n4684), .Z(n4682) );
  IV U2739 ( .A(n4685), .Z(n4683) );
  AN2 U2740 ( .A(U7_DATA1_53), .B(n4685), .Z(n4681) );
  OR2 U2741 ( .A(n4686), .B(n4687), .Z(n4685) );
  OR2 U2742 ( .A(n279), .B(n4688), .Z(n4687) );
  AN2 U2743 ( .A(ENCODER_DATA_IN[53]), .B(n4445), .Z(n4688) );
  AN2 U2744 ( .A(U15_Z_3), .B(n4446), .Z(n4686) );
  AN2 U2745 ( .A(n4689), .B(n4690), .Z(ENCODER_DATA_OUT[16]) );
  IV U2746 ( .A(n4691), .Z(n4690) );
  AN2 U2747 ( .A(n4692), .B(n4693), .Z(n4691) );
  OR2 U2748 ( .A(n4693), .B(n4692), .Z(n4689) );
  OR2 U2749 ( .A(n4694), .B(n4695), .Z(n4692) );
  AN2 U2750 ( .A(U7_DATA1_14), .B(n4696), .Z(n4695) );
  AN2 U2751 ( .A(U7_DATA1_33), .B(n4697), .Z(n4694) );
  IV U2752 ( .A(U7_DATA1_14), .Z(n4697) );
  OR2 U2753 ( .A(n4698), .B(n4699), .Z(n4693) );
  OR2 U2754 ( .A(n279), .B(n4700), .Z(n4699) );
  AN2 U2755 ( .A(ENCODER_DATA_IN[14]), .B(n4445), .Z(n4700) );
  AN2 U2756 ( .A(U34_Z_2), .B(n4446), .Z(n4698) );
  AN2 U2757 ( .A(TEST_PAT_SEED_A[47]), .B(n4391), .Z(n4675) );
  AN2 U2758 ( .A(TEST_PAT_SEED_B[47]), .B(n4392), .Z(n4673) );
  OR2 U2759 ( .A(n4701), .B(n4702), .Z(U5_Z_46) );
  OR2 U2760 ( .A(n4703), .B(n4704), .Z(n4702) );
  OR2 U2761 ( .A(n4705), .B(n4706), .Z(n4704) );
  AN2 U2762 ( .A(U7_DATA4_46), .B(n4384), .Z(n4706) );
  AN2 U2763 ( .A(U7_DATA6_46), .B(n4385), .Z(n4705) );
  AN2 U2764 ( .A(n2661), .B(U7_DATA1_46), .Z(n4703) );
  OR2 U2765 ( .A(n4707), .B(n4708), .Z(n4701) );
  OR2 U2766 ( .A(n4709), .B(n4710), .Z(n4708) );
  AN2 U2767 ( .A(n4390), .B(ENCODER_DATA_OUT[54]), .Z(n4710) );
  OR2 U2768 ( .A(n4711), .B(n4712), .Z(ENCODER_DATA_OUT[54]) );
  AN2 U2769 ( .A(n4713), .B(ENCODER_DATA_OUT[15]), .Z(n4712) );
  IV U2770 ( .A(n4714), .Z(n4711) );
  OR2 U2771 ( .A(ENCODER_DATA_OUT[15]), .B(n4713), .Z(n4714) );
  OR2 U2772 ( .A(n4715), .B(n4716), .Z(n4713) );
  AN2 U2773 ( .A(n4717), .B(n4718), .Z(n4716) );
  IV U2774 ( .A(n4719), .Z(n4717) );
  AN2 U2775 ( .A(U7_DATA1_52), .B(n4719), .Z(n4715) );
  OR2 U2776 ( .A(n4720), .B(n4721), .Z(n4719) );
  OR2 U2777 ( .A(n279), .B(n4722), .Z(n4721) );
  AN2 U2778 ( .A(ENCODER_DATA_IN[52]), .B(n4445), .Z(n4722) );
  AN2 U2779 ( .A(U15_Z_2), .B(n4446), .Z(n4720) );
  AN2 U2780 ( .A(n4723), .B(n4724), .Z(ENCODER_DATA_OUT[15]) );
  IV U2781 ( .A(n4725), .Z(n4724) );
  AN2 U2782 ( .A(n4726), .B(n4727), .Z(n4725) );
  OR2 U2783 ( .A(n4727), .B(n4726), .Z(n4723) );
  OR2 U2784 ( .A(n4728), .B(n4729), .Z(n4726) );
  AN2 U2785 ( .A(U7_DATA1_13), .B(n4730), .Z(n4729) );
  AN2 U2786 ( .A(U7_DATA1_32), .B(n4731), .Z(n4728) );
  IV U2787 ( .A(U7_DATA1_13), .Z(n4731) );
  OR2 U2788 ( .A(n4732), .B(n4733), .Z(n4727) );
  OR2 U2789 ( .A(n279), .B(n4734), .Z(n4733) );
  AN2 U2790 ( .A(ENCODER_DATA_IN[13]), .B(n4445), .Z(n4734) );
  AN2 U2791 ( .A(U34_Z_1), .B(n4446), .Z(n4732) );
  AN2 U2792 ( .A(TEST_PAT_SEED_A[46]), .B(n4391), .Z(n4709) );
  AN2 U2793 ( .A(TEST_PAT_SEED_B[46]), .B(n4392), .Z(n4707) );
  OR2 U2794 ( .A(n4735), .B(n4736), .Z(U5_Z_45) );
  OR2 U2795 ( .A(n4737), .B(n4738), .Z(n4736) );
  OR2 U2796 ( .A(n4739), .B(n4740), .Z(n4738) );
  AN2 U2797 ( .A(U7_DATA4_45), .B(n4384), .Z(n4740) );
  AN2 U2798 ( .A(U7_DATA6_45), .B(n4385), .Z(n4739) );
  AN2 U2799 ( .A(n2661), .B(U7_DATA1_45), .Z(n4737) );
  OR2 U2800 ( .A(n4741), .B(n4742), .Z(n4735) );
  OR2 U2801 ( .A(n4743), .B(n4744), .Z(n4742) );
  AN2 U2802 ( .A(n4390), .B(ENCODER_DATA_OUT[53]), .Z(n4744) );
  OR2 U2803 ( .A(n4745), .B(n4746), .Z(ENCODER_DATA_OUT[53]) );
  AN2 U2804 ( .A(n4747), .B(ENCODER_DATA_OUT[14]), .Z(n4746) );
  IV U2805 ( .A(n4748), .Z(n4745) );
  OR2 U2806 ( .A(ENCODER_DATA_OUT[14]), .B(n4747), .Z(n4748) );
  OR2 U2807 ( .A(n4749), .B(n4750), .Z(n4747) );
  AN2 U2808 ( .A(n4751), .B(n4752), .Z(n4750) );
  IV U2809 ( .A(n4753), .Z(n4751) );
  AN2 U2810 ( .A(U7_DATA1_51), .B(n4753), .Z(n4749) );
  OR2 U2811 ( .A(n4754), .B(n4755), .Z(n4753) );
  OR2 U2812 ( .A(n279), .B(n4756), .Z(n4755) );
  AN2 U2813 ( .A(ENCODER_DATA_IN[51]), .B(n4445), .Z(n4756) );
  AN2 U2814 ( .A(U15_Z_1), .B(n4446), .Z(n4754) );
  AN2 U2815 ( .A(n4757), .B(n4758), .Z(ENCODER_DATA_OUT[14]) );
  IV U2816 ( .A(n4759), .Z(n4758) );
  AN2 U2817 ( .A(n4760), .B(n4761), .Z(n4759) );
  OR2 U2818 ( .A(n4761), .B(n4760), .Z(n4757) );
  OR2 U2819 ( .A(n4762), .B(n4763), .Z(n4760) );
  AN2 U2820 ( .A(U7_DATA1_12), .B(n4764), .Z(n4763) );
  AN2 U2821 ( .A(U7_DATA1_31), .B(n4765), .Z(n4762) );
  IV U2822 ( .A(U7_DATA1_12), .Z(n4765) );
  OR2 U2823 ( .A(n4766), .B(n4767), .Z(n4761) );
  OR2 U2824 ( .A(n279), .B(n4768), .Z(n4767) );
  AN2 U2825 ( .A(ENCODER_DATA_IN[12]), .B(n4445), .Z(n4768) );
  AN2 U2826 ( .A(U33_Z_3), .B(n4446), .Z(n4766) );
  AN2 U2827 ( .A(TEST_PAT_SEED_A[45]), .B(n4391), .Z(n4743) );
  AN2 U2828 ( .A(TEST_PAT_SEED_B[45]), .B(n4392), .Z(n4741) );
  OR2 U2829 ( .A(n4769), .B(n4770), .Z(U5_Z_44) );
  OR2 U2830 ( .A(n4771), .B(n4772), .Z(n4770) );
  OR2 U2831 ( .A(n4773), .B(n4774), .Z(n4772) );
  AN2 U2832 ( .A(U7_DATA4_44), .B(n4384), .Z(n4774) );
  AN2 U2833 ( .A(U7_DATA6_44), .B(n4385), .Z(n4773) );
  AN2 U2834 ( .A(n2661), .B(U7_DATA1_44), .Z(n4771) );
  OR2 U2835 ( .A(n4775), .B(n4776), .Z(n4769) );
  OR2 U2836 ( .A(n4777), .B(n4778), .Z(n4776) );
  AN2 U2837 ( .A(n4390), .B(ENCODER_DATA_OUT[52]), .Z(n4778) );
  OR2 U2838 ( .A(n4779), .B(n4780), .Z(ENCODER_DATA_OUT[52]) );
  AN2 U2839 ( .A(n4781), .B(ENCODER_DATA_OUT[13]), .Z(n4780) );
  IV U2840 ( .A(n4782), .Z(n4779) );
  OR2 U2841 ( .A(ENCODER_DATA_OUT[13]), .B(n4781), .Z(n4782) );
  OR2 U2842 ( .A(n4783), .B(n4784), .Z(n4781) );
  AN2 U2843 ( .A(n4785), .B(n4786), .Z(n4784) );
  IV U2844 ( .A(n4787), .Z(n4785) );
  AN2 U2845 ( .A(U7_DATA1_50), .B(n4787), .Z(n4783) );
  OR2 U2846 ( .A(n4788), .B(n4789), .Z(n4787) );
  OR2 U2847 ( .A(n279), .B(n4790), .Z(n4789) );
  AN2 U2848 ( .A(ENCODER_DATA_IN[50]), .B(n4445), .Z(n4790) );
  AN2 U2849 ( .A(U15_Z_0), .B(n4446), .Z(n4788) );
  AN2 U2850 ( .A(n4791), .B(n4792), .Z(ENCODER_DATA_OUT[13]) );
  IV U2851 ( .A(n4793), .Z(n4792) );
  AN2 U2852 ( .A(n4794), .B(n4795), .Z(n4793) );
  OR2 U2853 ( .A(n4795), .B(n4794), .Z(n4791) );
  OR2 U2854 ( .A(n4796), .B(n4797), .Z(n4794) );
  AN2 U2855 ( .A(U7_DATA1_11), .B(n4798), .Z(n4797) );
  AN2 U2856 ( .A(U7_DATA1_30), .B(n4799), .Z(n4796) );
  IV U2857 ( .A(U7_DATA1_11), .Z(n4799) );
  OR2 U2858 ( .A(n4800), .B(n4801), .Z(n4795) );
  OR2 U2859 ( .A(n279), .B(n4802), .Z(n4801) );
  AN2 U2860 ( .A(ENCODER_DATA_IN[11]), .B(n4445), .Z(n4802) );
  AN2 U2861 ( .A(U33_Z_2), .B(n4446), .Z(n4800) );
  AN2 U2862 ( .A(TEST_PAT_SEED_A[44]), .B(n4391), .Z(n4777) );
  AN2 U2863 ( .A(TEST_PAT_SEED_B[44]), .B(n4392), .Z(n4775) );
  OR2 U2864 ( .A(n4803), .B(n4804), .Z(U5_Z_43) );
  OR2 U2865 ( .A(n4805), .B(n4806), .Z(n4804) );
  OR2 U2866 ( .A(n4807), .B(n4808), .Z(n4806) );
  AN2 U2867 ( .A(U7_DATA4_43), .B(n4384), .Z(n4808) );
  AN2 U2868 ( .A(U7_DATA6_43), .B(n4385), .Z(n4807) );
  AN2 U2869 ( .A(n2661), .B(U7_DATA1_43), .Z(n4805) );
  OR2 U2870 ( .A(n4809), .B(n4810), .Z(n4803) );
  OR2 U2871 ( .A(n4811), .B(n4812), .Z(n4810) );
  AN2 U2872 ( .A(n4390), .B(ENCODER_DATA_OUT[51]), .Z(n4812) );
  OR2 U2873 ( .A(n4813), .B(n4814), .Z(ENCODER_DATA_OUT[51]) );
  AN2 U2874 ( .A(n4815), .B(ENCODER_DATA_OUT[12]), .Z(n4814) );
  IV U2875 ( .A(n4816), .Z(n4813) );
  OR2 U2876 ( .A(ENCODER_DATA_OUT[12]), .B(n4815), .Z(n4816) );
  OR2 U2877 ( .A(n4817), .B(n4818), .Z(n4815) );
  AN2 U2878 ( .A(n4819), .B(n4820), .Z(n4818) );
  IV U2879 ( .A(n4821), .Z(n4819) );
  AN2 U2880 ( .A(U7_DATA1_49), .B(n4821), .Z(n4817) );
  OR2 U2881 ( .A(n4822), .B(n4823), .Z(n4821) );
  OR2 U2882 ( .A(n279), .B(n4824), .Z(n4823) );
  AN2 U2883 ( .A(ENCODER_DATA_IN[49]), .B(n4445), .Z(n4824) );
  AN2 U2884 ( .A(U16_Z_1), .B(n4446), .Z(n4822) );
  AN2 U2885 ( .A(TEST_PAT_SEED_A[43]), .B(n4391), .Z(n4811) );
  AN2 U2886 ( .A(TEST_PAT_SEED_B[43]), .B(n4392), .Z(n4809) );
  OR2 U2887 ( .A(n4825), .B(n4826), .Z(U5_Z_42) );
  OR2 U2888 ( .A(n4827), .B(n4828), .Z(n4826) );
  OR2 U2889 ( .A(n4829), .B(n4830), .Z(n4828) );
  AN2 U2890 ( .A(U7_DATA4_42), .B(n4384), .Z(n4830) );
  AN2 U2891 ( .A(U7_DATA6_42), .B(n4385), .Z(n4829) );
  AN2 U2892 ( .A(n2661), .B(U7_DATA1_42), .Z(n4827) );
  OR2 U2893 ( .A(n4831), .B(n4832), .Z(n4825) );
  OR2 U2894 ( .A(n4833), .B(n4834), .Z(n4832) );
  AN2 U2895 ( .A(n4390), .B(ENCODER_DATA_OUT[50]), .Z(n4834) );
  OR2 U2896 ( .A(n4835), .B(n4836), .Z(ENCODER_DATA_OUT[50]) );
  AN2 U2897 ( .A(n4837), .B(ENCODER_DATA_OUT[11]), .Z(n4836) );
  IV U2898 ( .A(n4838), .Z(n4835) );
  OR2 U2899 ( .A(ENCODER_DATA_OUT[11]), .B(n4837), .Z(n4838) );
  OR2 U2900 ( .A(n4839), .B(n4840), .Z(n4837) );
  AN2 U2901 ( .A(n4841), .B(n4842), .Z(n4840) );
  IV U2902 ( .A(n4843), .Z(n4841) );
  AN2 U2903 ( .A(U7_DATA1_48), .B(n4843), .Z(n4839) );
  OR2 U2904 ( .A(n4844), .B(n4845), .Z(n4843) );
  OR2 U2905 ( .A(n279), .B(n4846), .Z(n4845) );
  AN2 U2906 ( .A(ENCODER_DATA_IN[48]), .B(n4445), .Z(n4846) );
  AN2 U2907 ( .A(U16_Z_0), .B(n4446), .Z(n4844) );
  AN2 U2908 ( .A(TEST_PAT_SEED_A[42]), .B(n4391), .Z(n4833) );
  AN2 U2909 ( .A(TEST_PAT_SEED_B[42]), .B(n4392), .Z(n4831) );
  OR2 U2910 ( .A(n4847), .B(n4848), .Z(U5_Z_41) );
  OR2 U2911 ( .A(n4849), .B(n4850), .Z(n4848) );
  OR2 U2912 ( .A(n4851), .B(n4852), .Z(n4850) );
  AN2 U2913 ( .A(U7_DATA4_41), .B(n4384), .Z(n4852) );
  AN2 U2914 ( .A(U7_DATA6_41), .B(n4385), .Z(n4851) );
  AN2 U2915 ( .A(n2661), .B(U7_DATA1_41), .Z(n4849) );
  OR2 U2916 ( .A(n4853), .B(n4854), .Z(n4847) );
  OR2 U2917 ( .A(n4855), .B(n4856), .Z(n4854) );
  AN2 U2918 ( .A(n4390), .B(ENCODER_DATA_OUT[49]), .Z(n4856) );
  OR2 U2919 ( .A(n4857), .B(n4858), .Z(ENCODER_DATA_OUT[49]) );
  AN2 U2920 ( .A(n4859), .B(ENCODER_DATA_OUT[10]), .Z(n4858) );
  IV U2921 ( .A(n4860), .Z(n4857) );
  OR2 U2922 ( .A(ENCODER_DATA_OUT[10]), .B(n4859), .Z(n4860) );
  OR2 U2923 ( .A(n4861), .B(n4862), .Z(n4859) );
  AN2 U2924 ( .A(n4863), .B(n4864), .Z(n4862) );
  IV U2925 ( .A(n4865), .Z(n4863) );
  AN2 U2926 ( .A(U7_DATA1_47), .B(n4865), .Z(n4861) );
  OR2 U2927 ( .A(n4866), .B(n4867), .Z(n4865) );
  OR2 U2928 ( .A(n279), .B(n4868), .Z(n4867) );
  AN2 U2929 ( .A(ENCODER_DATA_IN[47]), .B(n4445), .Z(n4868) );
  AN2 U2930 ( .A(U17_Z_4), .B(n4446), .Z(n4866) );
  AN2 U2931 ( .A(TEST_PAT_SEED_A[41]), .B(n4391), .Z(n4855) );
  AN2 U2932 ( .A(TEST_PAT_SEED_B[41]), .B(n4392), .Z(n4853) );
  OR2 U2933 ( .A(n4869), .B(n4870), .Z(U5_Z_40) );
  OR2 U2934 ( .A(n4871), .B(n4872), .Z(n4870) );
  OR2 U2935 ( .A(n4873), .B(n4874), .Z(n4872) );
  AN2 U2936 ( .A(U7_DATA4_40), .B(n4384), .Z(n4874) );
  AN2 U2937 ( .A(U7_DATA6_40), .B(n4385), .Z(n4873) );
  AN2 U2938 ( .A(n2661), .B(U7_DATA1_40), .Z(n4871) );
  OR2 U2939 ( .A(n4875), .B(n4876), .Z(n4869) );
  OR2 U2940 ( .A(n4877), .B(n4878), .Z(n4876) );
  AN2 U2941 ( .A(n4390), .B(ENCODER_DATA_OUT[48]), .Z(n4878) );
  OR2 U2942 ( .A(n4879), .B(n4880), .Z(ENCODER_DATA_OUT[48]) );
  AN2 U2943 ( .A(n4881), .B(ENCODER_DATA_OUT[9]), .Z(n4880) );
  IV U2944 ( .A(n4882), .Z(n4879) );
  OR2 U2945 ( .A(ENCODER_DATA_OUT[9]), .B(n4881), .Z(n4882) );
  OR2 U2946 ( .A(n4883), .B(n4884), .Z(n4881) );
  AN2 U2947 ( .A(n4885), .B(n4886), .Z(n4884) );
  IV U2948 ( .A(n4887), .Z(n4885) );
  AN2 U2949 ( .A(U7_DATA1_46), .B(n4887), .Z(n4883) );
  OR2 U2950 ( .A(n4888), .B(n4889), .Z(n4887) );
  OR2 U2951 ( .A(n279), .B(n4890), .Z(n4889) );
  AN2 U2952 ( .A(ENCODER_DATA_IN[46]), .B(n4445), .Z(n4890) );
  AN2 U2953 ( .A(U17_Z_3), .B(n4446), .Z(n4888) );
  AN2 U2954 ( .A(TEST_PAT_SEED_A[40]), .B(n4391), .Z(n4877) );
  AN2 U2955 ( .A(TEST_PAT_SEED_B[40]), .B(n4392), .Z(n4875) );
  OR2 U2956 ( .A(n4891), .B(n4892), .Z(U5_Z_4) );
  OR2 U2957 ( .A(n4893), .B(n4894), .Z(n4892) );
  OR2 U2958 ( .A(n4895), .B(n4896), .Z(n4894) );
  AN2 U2959 ( .A(U7_DATA4_4), .B(n4384), .Z(n4896) );
  AN2 U2960 ( .A(U7_DATA6_4), .B(n4385), .Z(n4895) );
  AN2 U2961 ( .A(n2661), .B(U7_DATA1_4), .Z(n4893) );
  OR2 U2962 ( .A(n4897), .B(n4898), .Z(n4891) );
  OR2 U2963 ( .A(n4899), .B(n4900), .Z(n4898) );
  AN2 U2964 ( .A(n4390), .B(ENCODER_DATA_OUT[12]), .Z(n4900) );
  AN2 U2965 ( .A(n4901), .B(n4902), .Z(ENCODER_DATA_OUT[12]) );
  IV U2966 ( .A(n4903), .Z(n4902) );
  AN2 U2967 ( .A(n4904), .B(n4905), .Z(n4903) );
  OR2 U2968 ( .A(n4905), .B(n4904), .Z(n4901) );
  OR2 U2969 ( .A(n4906), .B(n4907), .Z(n4904) );
  AN2 U2970 ( .A(U7_DATA1_10), .B(n4908), .Z(n4907) );
  AN2 U2971 ( .A(U7_DATA1_29), .B(n4909), .Z(n4906) );
  IV U2972 ( .A(U7_DATA1_10), .Z(n4909) );
  OR2 U2973 ( .A(n4910), .B(n4911), .Z(n4905) );
  OR2 U2974 ( .A(n279), .B(n4912), .Z(n4911) );
  AN2 U2975 ( .A(ENCODER_DATA_IN[10]), .B(n4445), .Z(n4912) );
  AN2 U2976 ( .A(U33_Z_1), .B(n4446), .Z(n4910) );
  AN2 U2977 ( .A(TEST_PAT_SEED_A[4]), .B(n4391), .Z(n4899) );
  AN2 U2978 ( .A(TEST_PAT_SEED_B[4]), .B(n4392), .Z(n4897) );
  OR2 U2979 ( .A(n4913), .B(n4914), .Z(U5_Z_39) );
  OR2 U2980 ( .A(n4915), .B(n4916), .Z(n4914) );
  OR2 U2981 ( .A(n4917), .B(n4918), .Z(n4916) );
  AN2 U2982 ( .A(U7_DATA4_39), .B(n4384), .Z(n4918) );
  AN2 U2983 ( .A(U7_DATA6_39), .B(n4385), .Z(n4917) );
  AN2 U2984 ( .A(n2661), .B(U7_DATA1_39), .Z(n4915) );
  OR2 U2985 ( .A(n4919), .B(n4920), .Z(n4913) );
  OR2 U2986 ( .A(n4921), .B(n4922), .Z(n4920) );
  AN2 U2987 ( .A(n4390), .B(ENCODER_DATA_OUT[47]), .Z(n4922) );
  OR2 U2988 ( .A(n4923), .B(n4924), .Z(ENCODER_DATA_OUT[47]) );
  AN2 U2989 ( .A(n4925), .B(ENCODER_DATA_OUT[8]), .Z(n4924) );
  IV U2990 ( .A(n4926), .Z(n4923) );
  OR2 U2991 ( .A(ENCODER_DATA_OUT[8]), .B(n4925), .Z(n4926) );
  OR2 U2992 ( .A(n4927), .B(n4928), .Z(n4925) );
  AN2 U2993 ( .A(n4929), .B(n4930), .Z(n4928) );
  IV U2994 ( .A(n4931), .Z(n4929) );
  AN2 U2995 ( .A(U7_DATA1_45), .B(n4931), .Z(n4927) );
  OR2 U2996 ( .A(n4932), .B(n4933), .Z(n4931) );
  OR2 U2997 ( .A(n279), .B(n4934), .Z(n4933) );
  AN2 U2998 ( .A(ENCODER_DATA_IN[45]), .B(n4445), .Z(n4934) );
  AN2 U2999 ( .A(U17_Z_2), .B(n4446), .Z(n4932) );
  AN2 U3000 ( .A(TEST_PAT_SEED_A[39]), .B(n4391), .Z(n4921) );
  AN2 U3001 ( .A(TEST_PAT_SEED_B[39]), .B(n4392), .Z(n4919) );
  OR2 U3002 ( .A(n4935), .B(n4936), .Z(U5_Z_38) );
  OR2 U3003 ( .A(n4937), .B(n4938), .Z(n4936) );
  OR2 U3004 ( .A(n4939), .B(n4940), .Z(n4938) );
  AN2 U3005 ( .A(U7_DATA4_38), .B(n4384), .Z(n4940) );
  AN2 U3006 ( .A(U7_DATA6_38), .B(n4385), .Z(n4939) );
  AN2 U3007 ( .A(n2661), .B(U7_DATA1_38), .Z(n4937) );
  OR2 U3008 ( .A(n4941), .B(n4942), .Z(n4935) );
  OR2 U3009 ( .A(n4943), .B(n4944), .Z(n4942) );
  AN2 U3010 ( .A(n4390), .B(ENCODER_DATA_OUT[46]), .Z(n4944) );
  OR2 U3011 ( .A(n4945), .B(n4946), .Z(ENCODER_DATA_OUT[46]) );
  AN2 U3012 ( .A(n4947), .B(ENCODER_DATA_OUT[7]), .Z(n4946) );
  IV U3013 ( .A(n4948), .Z(n4945) );
  OR2 U3014 ( .A(ENCODER_DATA_OUT[7]), .B(n4947), .Z(n4948) );
  OR2 U3015 ( .A(n4949), .B(n4950), .Z(n4947) );
  AN2 U3016 ( .A(n4951), .B(n4952), .Z(n4950) );
  IV U3017 ( .A(n4953), .Z(n4951) );
  AN2 U3018 ( .A(U7_DATA1_44), .B(n4953), .Z(n4949) );
  OR2 U3019 ( .A(n4954), .B(n4955), .Z(n4953) );
  OR2 U3020 ( .A(n279), .B(n4956), .Z(n4955) );
  AN2 U3021 ( .A(ENCODER_DATA_IN[44]), .B(n4445), .Z(n4956) );
  AN2 U3022 ( .A(U17_Z_1), .B(n4446), .Z(n4954) );
  AN2 U3023 ( .A(TEST_PAT_SEED_A[38]), .B(n4391), .Z(n4943) );
  AN2 U3024 ( .A(TEST_PAT_SEED_B[38]), .B(n4392), .Z(n4941) );
  OR2 U3025 ( .A(n4957), .B(n4958), .Z(U5_Z_37) );
  OR2 U3026 ( .A(n4959), .B(n4960), .Z(n4958) );
  OR2 U3027 ( .A(n4961), .B(n4962), .Z(n4960) );
  AN2 U3028 ( .A(U7_DATA4_37), .B(n4384), .Z(n4962) );
  AN2 U3029 ( .A(U7_DATA6_37), .B(n4385), .Z(n4961) );
  AN2 U3030 ( .A(n2661), .B(U7_DATA1_37), .Z(n4959) );
  OR2 U3031 ( .A(n4963), .B(n4964), .Z(n4957) );
  OR2 U3032 ( .A(n4965), .B(n4966), .Z(n4964) );
  AN2 U3033 ( .A(n4390), .B(ENCODER_DATA_OUT[45]), .Z(n4966) );
  OR2 U3034 ( .A(n4967), .B(n4968), .Z(ENCODER_DATA_OUT[45]) );
  AN2 U3035 ( .A(n4969), .B(ENCODER_DATA_OUT[6]), .Z(n4968) );
  IV U3036 ( .A(n4970), .Z(n4967) );
  OR2 U3037 ( .A(ENCODER_DATA_OUT[6]), .B(n4969), .Z(n4970) );
  OR2 U3038 ( .A(n4971), .B(n4972), .Z(n4969) );
  IV U3039 ( .A(n4973), .Z(n4972) );
  OR2 U3040 ( .A(n4974), .B(U7_DATA1_43), .Z(n4973) );
  AN2 U3041 ( .A(U7_DATA1_43), .B(n4974), .Z(n4971) );
  OR2 U3042 ( .A(n4975), .B(n4976), .Z(n4974) );
  OR2 U3043 ( .A(n279), .B(n4977), .Z(n4976) );
  AN2 U3044 ( .A(ENCODER_DATA_IN[43]), .B(n4445), .Z(n4977) );
  AN2 U3045 ( .A(U17_Z_0), .B(n4446), .Z(n4975) );
  AN2 U3046 ( .A(TEST_PAT_SEED_A[37]), .B(n4391), .Z(n4965) );
  AN2 U3047 ( .A(TEST_PAT_SEED_B[37]), .B(n4392), .Z(n4963) );
  OR2 U3048 ( .A(n4978), .B(n4979), .Z(U5_Z_36) );
  OR2 U3049 ( .A(n4980), .B(n4981), .Z(n4979) );
  OR2 U3050 ( .A(n4982), .B(n4983), .Z(n4981) );
  AN2 U3051 ( .A(U7_DATA4_36), .B(n4384), .Z(n4983) );
  AN2 U3052 ( .A(U7_DATA6_36), .B(n4385), .Z(n4982) );
  AN2 U3053 ( .A(n2661), .B(U7_DATA1_36), .Z(n4980) );
  OR2 U3054 ( .A(n4984), .B(n4985), .Z(n4978) );
  OR2 U3055 ( .A(n4986), .B(n4987), .Z(n4985) );
  AN2 U3056 ( .A(n4390), .B(ENCODER_DATA_OUT[44]), .Z(n4987) );
  OR2 U3057 ( .A(n4988), .B(n4989), .Z(ENCODER_DATA_OUT[44]) );
  AN2 U3058 ( .A(n4990), .B(ENCODER_DATA_OUT[5]), .Z(n4989) );
  IV U3059 ( .A(n4991), .Z(n4988) );
  OR2 U3060 ( .A(ENCODER_DATA_OUT[5]), .B(n4990), .Z(n4991) );
  OR2 U3061 ( .A(n4992), .B(n4993), .Z(n4990) );
  IV U3062 ( .A(n4994), .Z(n4993) );
  OR2 U3063 ( .A(n4995), .B(U7_DATA1_42), .Z(n4994) );
  AN2 U3064 ( .A(U7_DATA1_42), .B(n4995), .Z(n4992) );
  OR2 U3065 ( .A(n4996), .B(n4997), .Z(n4995) );
  OR2 U3066 ( .A(n279), .B(n4998), .Z(n4997) );
  AN2 U3067 ( .A(ENCODER_DATA_IN[42]), .B(n4445), .Z(n4998) );
  AN2 U3068 ( .A(U18_Z_1), .B(n4446), .Z(n4996) );
  AN2 U3069 ( .A(TEST_PAT_SEED_A[36]), .B(n4391), .Z(n4986) );
  AN2 U3070 ( .A(TEST_PAT_SEED_B[36]), .B(n4392), .Z(n4984) );
  OR2 U3071 ( .A(n4999), .B(n5000), .Z(U5_Z_35) );
  OR2 U3072 ( .A(n5001), .B(n5002), .Z(n5000) );
  OR2 U3073 ( .A(n5003), .B(n5004), .Z(n5002) );
  AN2 U3074 ( .A(U7_DATA4_35), .B(n4384), .Z(n5004) );
  AN2 U3075 ( .A(U7_DATA6_35), .B(n4385), .Z(n5003) );
  AN2 U3076 ( .A(n2661), .B(U7_DATA1_35), .Z(n5001) );
  OR2 U3077 ( .A(n5005), .B(n5006), .Z(n4999) );
  OR2 U3078 ( .A(n5007), .B(n5008), .Z(n5006) );
  AN2 U3079 ( .A(n4390), .B(ENCODER_DATA_OUT[43]), .Z(n5008) );
  OR2 U3080 ( .A(n5009), .B(n5010), .Z(ENCODER_DATA_OUT[43]) );
  AN2 U3081 ( .A(n5011), .B(ENCODER_DATA_OUT[4]), .Z(n5010) );
  IV U3082 ( .A(n5012), .Z(n5009) );
  OR2 U3083 ( .A(ENCODER_DATA_OUT[4]), .B(n5011), .Z(n5012) );
  OR2 U3084 ( .A(n5013), .B(n5014), .Z(n5011) );
  IV U3085 ( .A(n5015), .Z(n5014) );
  OR2 U3086 ( .A(n5016), .B(U7_DATA1_41), .Z(n5015) );
  AN2 U3087 ( .A(U7_DATA1_41), .B(n5016), .Z(n5013) );
  OR2 U3088 ( .A(n5017), .B(n5018), .Z(n5016) );
  OR2 U3089 ( .A(n279), .B(n5019), .Z(n5018) );
  AN2 U3090 ( .A(ENCODER_DATA_IN[41]), .B(n4445), .Z(n5019) );
  AN2 U3091 ( .A(U18_Z_0), .B(n4446), .Z(n5017) );
  AN2 U3092 ( .A(TEST_PAT_SEED_A[35]), .B(n4391), .Z(n5007) );
  AN2 U3093 ( .A(TEST_PAT_SEED_B[35]), .B(n4392), .Z(n5005) );
  OR2 U3094 ( .A(n5020), .B(n5021), .Z(U5_Z_34) );
  OR2 U3095 ( .A(n5022), .B(n5023), .Z(n5021) );
  OR2 U3096 ( .A(n5024), .B(n5025), .Z(n5023) );
  AN2 U3097 ( .A(U7_DATA4_34), .B(n4384), .Z(n5025) );
  AN2 U3098 ( .A(U7_DATA6_34), .B(n4385), .Z(n5024) );
  AN2 U3099 ( .A(n2661), .B(U7_DATA1_34), .Z(n5022) );
  OR2 U3100 ( .A(n5026), .B(n5027), .Z(n5020) );
  OR2 U3101 ( .A(n5028), .B(n5029), .Z(n5027) );
  AN2 U3102 ( .A(n4390), .B(ENCODER_DATA_OUT[42]), .Z(n5029) );
  OR2 U3103 ( .A(n5030), .B(n5031), .Z(ENCODER_DATA_OUT[42]) );
  AN2 U3104 ( .A(n5032), .B(ENCODER_DATA_OUT[3]), .Z(n5031) );
  IV U3105 ( .A(n5033), .Z(n5030) );
  OR2 U3106 ( .A(ENCODER_DATA_OUT[3]), .B(n5032), .Z(n5033) );
  OR2 U3107 ( .A(n5034), .B(n5035), .Z(n5032) );
  IV U3108 ( .A(n5036), .Z(n5035) );
  OR2 U3109 ( .A(n5037), .B(U7_DATA1_40), .Z(n5036) );
  AN2 U3110 ( .A(U7_DATA1_40), .B(n5037), .Z(n5034) );
  OR2 U3111 ( .A(n5038), .B(n5039), .Z(n5037) );
  OR2 U3112 ( .A(n279), .B(n5040), .Z(n5039) );
  AN2 U3113 ( .A(ENCODER_DATA_IN[40]), .B(n4445), .Z(n5040) );
  AN2 U3114 ( .A(U19_Z_0), .B(n4446), .Z(n5038) );
  AN2 U3115 ( .A(TEST_PAT_SEED_A[34]), .B(n4391), .Z(n5028) );
  AN2 U3116 ( .A(TEST_PAT_SEED_B[34]), .B(n4392), .Z(n5026) );
  OR2 U3117 ( .A(n5041), .B(n5042), .Z(U5_Z_33) );
  OR2 U3118 ( .A(n5043), .B(n5044), .Z(n5042) );
  OR2 U3119 ( .A(n5045), .B(n5046), .Z(n5044) );
  AN2 U3120 ( .A(U7_DATA4_33), .B(n4384), .Z(n5046) );
  AN2 U3121 ( .A(U7_DATA6_33), .B(n4385), .Z(n5045) );
  AN2 U3122 ( .A(n2661), .B(U7_DATA1_33), .Z(n5043) );
  OR2 U3123 ( .A(n5047), .B(n5048), .Z(n5041) );
  OR2 U3124 ( .A(n5049), .B(n5050), .Z(n5048) );
  AN2 U3125 ( .A(n4390), .B(ENCODER_DATA_OUT[41]), .Z(n5050) );
  OR2 U3126 ( .A(n5051), .B(n5052), .Z(ENCODER_DATA_OUT[41]) );
  AN2 U3127 ( .A(n5053), .B(ENCODER_DATA_OUT[2]), .Z(n5052) );
  IV U3128 ( .A(n5054), .Z(n5051) );
  OR2 U3129 ( .A(ENCODER_DATA_OUT[2]), .B(n5053), .Z(n5054) );
  OR2 U3130 ( .A(n5055), .B(n5056), .Z(n5053) );
  IV U3131 ( .A(n5057), .Z(n5056) );
  OR2 U3132 ( .A(n5058), .B(U7_DATA1_39), .Z(n5057) );
  AN2 U3133 ( .A(U7_DATA1_39), .B(n5058), .Z(n5055) );
  OR2 U3134 ( .A(n5059), .B(n5060), .Z(n5058) );
  OR2 U3135 ( .A(n279), .B(n5061), .Z(n5060) );
  AN2 U3136 ( .A(ENCODER_DATA_IN[39]), .B(n4445), .Z(n5061) );
  AN2 U3137 ( .A(U20_Z_2), .B(n4446), .Z(n5059) );
  AN2 U3138 ( .A(TEST_PAT_SEED_A[33]), .B(n4391), .Z(n5049) );
  AN2 U3139 ( .A(TEST_PAT_SEED_B[33]), .B(n4392), .Z(n5047) );
  OR2 U3140 ( .A(n5062), .B(n5063), .Z(U5_Z_32) );
  OR2 U3141 ( .A(n5064), .B(n5065), .Z(n5063) );
  OR2 U3142 ( .A(n5066), .B(n5067), .Z(n5065) );
  AN2 U3143 ( .A(U7_DATA4_32), .B(n4384), .Z(n5067) );
  AN2 U3144 ( .A(U7_DATA6_32), .B(n4385), .Z(n5066) );
  AN2 U3145 ( .A(n2661), .B(U7_DATA1_32), .Z(n5064) );
  OR2 U3146 ( .A(n5068), .B(n5069), .Z(n5062) );
  OR2 U3147 ( .A(n5070), .B(n5071), .Z(n5069) );
  AN2 U3148 ( .A(ENCODER_DATA_OUT[40]), .B(n4390), .Z(n5071) );
  IV U3149 ( .A(n5072), .Z(ENCODER_DATA_OUT[40]) );
  OR2 U3150 ( .A(n5073), .B(n5074), .Z(n5072) );
  AN2 U3151 ( .A(n5075), .B(n5076), .Z(n5074) );
  AN2 U3152 ( .A(n5077), .B(n5078), .Z(n5076) );
  OR2 U3153 ( .A(U7_DATA1_38), .B(n4574), .Z(n5078) );
  OR2 U3154 ( .A(U7_DATA1_57), .B(n5079), .Z(n5077) );
  IV U3155 ( .A(n5080), .Z(n5075) );
  AN2 U3156 ( .A(n5081), .B(n5080), .Z(n5073) );
  OR2 U3157 ( .A(n5082), .B(n5083), .Z(n5080) );
  OR2 U3158 ( .A(n279), .B(n5084), .Z(n5083) );
  AN2 U3159 ( .A(ENCODER_DATA_IN[38]), .B(n4445), .Z(n5084) );
  AN2 U3160 ( .A(U20_Z_1), .B(n4446), .Z(n5082) );
  OR2 U3161 ( .A(n5085), .B(n5086), .Z(n5081) );
  AN2 U3162 ( .A(U7_DATA1_38), .B(n4574), .Z(n5086) );
  IV U3163 ( .A(U7_DATA1_57), .Z(n4574) );
  AN2 U3164 ( .A(U7_DATA1_57), .B(n5079), .Z(n5085) );
  AN2 U3165 ( .A(TEST_PAT_SEED_A[32]), .B(n4391), .Z(n5070) );
  AN2 U3166 ( .A(TEST_PAT_SEED_B[32]), .B(n4392), .Z(n5068) );
  OR2 U3167 ( .A(n5087), .B(n5088), .Z(U5_Z_31) );
  OR2 U3168 ( .A(n5089), .B(n5090), .Z(n5088) );
  OR2 U3169 ( .A(n5091), .B(n5092), .Z(n5090) );
  AN2 U3170 ( .A(U7_DATA4_31), .B(n4384), .Z(n5092) );
  AN2 U3171 ( .A(U7_DATA6_31), .B(n4385), .Z(n5091) );
  AN2 U3172 ( .A(n2661), .B(U7_DATA1_31), .Z(n5089) );
  OR2 U3173 ( .A(n5093), .B(n5094), .Z(n5087) );
  OR2 U3174 ( .A(n5095), .B(n5096), .Z(n5094) );
  AN2 U3175 ( .A(ENCODER_DATA_OUT[39]), .B(n4390), .Z(n5096) );
  IV U3176 ( .A(n5097), .Z(ENCODER_DATA_OUT[39]) );
  OR2 U3177 ( .A(n5098), .B(n5099), .Z(n5097) );
  AN2 U3178 ( .A(n5100), .B(n5101), .Z(n5099) );
  AN2 U3179 ( .A(n5102), .B(n5103), .Z(n5101) );
  OR2 U3180 ( .A(U7_DATA1_37), .B(n4596), .Z(n5103) );
  OR2 U3181 ( .A(U7_DATA1_56), .B(n5104), .Z(n5102) );
  IV U3182 ( .A(n5105), .Z(n5100) );
  AN2 U3183 ( .A(n5106), .B(n5105), .Z(n5098) );
  OR2 U3184 ( .A(n5107), .B(n5108), .Z(n5105) );
  OR2 U3185 ( .A(n279), .B(n5109), .Z(n5108) );
  AN2 U3186 ( .A(ENCODER_DATA_IN[37]), .B(n4445), .Z(n5109) );
  AN2 U3187 ( .A(U20_Z_0), .B(n4446), .Z(n5107) );
  OR2 U3188 ( .A(n5110), .B(n5111), .Z(n5106) );
  AN2 U3189 ( .A(U7_DATA1_37), .B(n4596), .Z(n5111) );
  IV U3190 ( .A(U7_DATA1_56), .Z(n4596) );
  AN2 U3191 ( .A(U7_DATA1_56), .B(n5104), .Z(n5110) );
  AN2 U3192 ( .A(TEST_PAT_SEED_A[31]), .B(n4391), .Z(n5095) );
  AN2 U3193 ( .A(TEST_PAT_SEED_B[31]), .B(n4392), .Z(n5093) );
  OR2 U3194 ( .A(n5112), .B(n5113), .Z(U5_Z_30) );
  OR2 U3195 ( .A(n5114), .B(n5115), .Z(n5113) );
  OR2 U3196 ( .A(n5116), .B(n5117), .Z(n5115) );
  AN2 U3197 ( .A(U7_DATA4_30), .B(n4384), .Z(n5117) );
  AN2 U3198 ( .A(U7_DATA6_30), .B(n4385), .Z(n5116) );
  AN2 U3199 ( .A(n2661), .B(U7_DATA1_30), .Z(n5114) );
  OR2 U3200 ( .A(n5118), .B(n5119), .Z(n5112) );
  OR2 U3201 ( .A(n5120), .B(n5121), .Z(n5119) );
  AN2 U3202 ( .A(ENCODER_DATA_OUT[38]), .B(n4390), .Z(n5121) );
  IV U3203 ( .A(n5122), .Z(ENCODER_DATA_OUT[38]) );
  OR2 U3204 ( .A(n5123), .B(n5124), .Z(n5122) );
  AN2 U3205 ( .A(n5125), .B(n5126), .Z(n5124) );
  AN2 U3206 ( .A(n5127), .B(n5128), .Z(n5126) );
  OR2 U3207 ( .A(U7_DATA1_36), .B(n4628), .Z(n5128) );
  OR2 U3208 ( .A(U7_DATA1_55), .B(n5129), .Z(n5127) );
  IV U3209 ( .A(n5130), .Z(n5125) );
  AN2 U3210 ( .A(n5131), .B(n5130), .Z(n5123) );
  OR2 U3211 ( .A(n5132), .B(n5133), .Z(n5130) );
  OR2 U3212 ( .A(n279), .B(n5134), .Z(n5133) );
  AN2 U3213 ( .A(ENCODER_DATA_IN[36]), .B(n4445), .Z(n5134) );
  AN2 U3214 ( .A(U23_Z_0), .B(n4446), .Z(n5132) );
  OR2 U3215 ( .A(n5135), .B(n5136), .Z(n5131) );
  AN2 U3216 ( .A(U7_DATA1_36), .B(n4628), .Z(n5136) );
  IV U3217 ( .A(U7_DATA1_55), .Z(n4628) );
  AN2 U3218 ( .A(U7_DATA1_55), .B(n5129), .Z(n5135) );
  AN2 U3219 ( .A(TEST_PAT_SEED_A[30]), .B(n4391), .Z(n5120) );
  AN2 U3220 ( .A(TEST_PAT_SEED_B[30]), .B(n4392), .Z(n5118) );
  OR2 U3221 ( .A(n5137), .B(n5138), .Z(U5_Z_3) );
  OR2 U3222 ( .A(n5139), .B(n5140), .Z(n5138) );
  OR2 U3223 ( .A(n5141), .B(n5142), .Z(n5140) );
  AN2 U3224 ( .A(U7_DATA4_3), .B(n4384), .Z(n5142) );
  AN2 U3225 ( .A(U7_DATA6_3), .B(n4385), .Z(n5141) );
  AN2 U3226 ( .A(n2661), .B(U7_DATA1_3), .Z(n5139) );
  OR2 U3227 ( .A(n5143), .B(n5144), .Z(n5137) );
  OR2 U3228 ( .A(n5145), .B(n5146), .Z(n5144) );
  AN2 U3229 ( .A(n4390), .B(ENCODER_DATA_OUT[11]), .Z(n5146) );
  AN2 U3230 ( .A(n5147), .B(n5148), .Z(ENCODER_DATA_OUT[11]) );
  IV U3231 ( .A(n5149), .Z(n5148) );
  AN2 U3232 ( .A(n5150), .B(n5151), .Z(n5149) );
  OR2 U3233 ( .A(n5151), .B(n5150), .Z(n5147) );
  OR2 U3234 ( .A(n5152), .B(n5153), .Z(n5150) );
  AN2 U3235 ( .A(U7_DATA1_28), .B(n5154), .Z(n5153) );
  IV U3236 ( .A(U7_DATA1_9), .Z(n5154) );
  AN2 U3237 ( .A(U7_DATA1_9), .B(n5155), .Z(n5152) );
  OR2 U3238 ( .A(n5156), .B(n5157), .Z(n5151) );
  OR2 U3239 ( .A(n279), .B(n5158), .Z(n5157) );
  AN2 U3240 ( .A(ENCODER_DATA_IN[9]), .B(n4445), .Z(n5158) );
  AN2 U3241 ( .A(U33_Z_0), .B(n4446), .Z(n5156) );
  AN2 U3242 ( .A(TEST_PAT_SEED_A[3]), .B(n4391), .Z(n5145) );
  AN2 U3243 ( .A(TEST_PAT_SEED_B[3]), .B(n4392), .Z(n5143) );
  OR2 U3244 ( .A(n5159), .B(n5160), .Z(U5_Z_29) );
  OR2 U3245 ( .A(n5161), .B(n5162), .Z(n5160) );
  OR2 U3246 ( .A(n5163), .B(n5164), .Z(n5162) );
  AN2 U3247 ( .A(U7_DATA4_29), .B(n4384), .Z(n5164) );
  AN2 U3248 ( .A(U7_DATA6_29), .B(n4385), .Z(n5163) );
  AN2 U3249 ( .A(n2661), .B(U7_DATA1_29), .Z(n5161) );
  OR2 U3250 ( .A(n5165), .B(n5166), .Z(n5159) );
  OR2 U3251 ( .A(n5167), .B(n5168), .Z(n5166) );
  AN2 U3252 ( .A(ENCODER_DATA_OUT[37]), .B(n4390), .Z(n5168) );
  IV U3253 ( .A(n5169), .Z(ENCODER_DATA_OUT[37]) );
  OR2 U3254 ( .A(n5170), .B(n5171), .Z(n5169) );
  AN2 U3255 ( .A(n5172), .B(n5173), .Z(n5171) );
  AN2 U3256 ( .A(n5174), .B(n5175), .Z(n5173) );
  OR2 U3257 ( .A(U7_DATA1_35), .B(n4650), .Z(n5175) );
  OR2 U3258 ( .A(U7_DATA1_54), .B(n5176), .Z(n5174) );
  IV U3259 ( .A(n5177), .Z(n5172) );
  AN2 U3260 ( .A(n5178), .B(n5177), .Z(n5170) );
  OR2 U3261 ( .A(n5179), .B(n5180), .Z(n5177) );
  OR2 U3262 ( .A(n279), .B(n5181), .Z(n5180) );
  AN2 U3263 ( .A(ENCODER_DATA_IN[35]), .B(n4445), .Z(n5181) );
  AN2 U3264 ( .A(U24_Z_1), .B(n4446), .Z(n5179) );
  OR2 U3265 ( .A(n5182), .B(n5183), .Z(n5178) );
  AN2 U3266 ( .A(U7_DATA1_35), .B(n4650), .Z(n5183) );
  IV U3267 ( .A(U7_DATA1_54), .Z(n4650) );
  AN2 U3268 ( .A(U7_DATA1_54), .B(n5176), .Z(n5182) );
  AN2 U3269 ( .A(TEST_PAT_SEED_A[29]), .B(n4391), .Z(n5167) );
  AN2 U3270 ( .A(TEST_PAT_SEED_B[29]), .B(n4392), .Z(n5165) );
  OR2 U3271 ( .A(n5184), .B(n5185), .Z(U5_Z_28) );
  OR2 U3272 ( .A(n5186), .B(n5187), .Z(n5185) );
  OR2 U3273 ( .A(n5188), .B(n5189), .Z(n5187) );
  AN2 U3274 ( .A(U7_DATA4_28), .B(n4384), .Z(n5189) );
  AN2 U3275 ( .A(U7_DATA6_28), .B(n4385), .Z(n5188) );
  AN2 U3276 ( .A(n2661), .B(U7_DATA1_28), .Z(n5186) );
  OR2 U3277 ( .A(n5190), .B(n5191), .Z(n5184) );
  OR2 U3278 ( .A(n5192), .B(n5193), .Z(n5191) );
  AN2 U3279 ( .A(ENCODER_DATA_OUT[36]), .B(n4390), .Z(n5193) );
  IV U3280 ( .A(n5194), .Z(ENCODER_DATA_OUT[36]) );
  OR2 U3281 ( .A(n5195), .B(n5196), .Z(n5194) );
  AN2 U3282 ( .A(n5197), .B(n5198), .Z(n5196) );
  AN2 U3283 ( .A(n5199), .B(n5200), .Z(n5198) );
  OR2 U3284 ( .A(U7_DATA1_34), .B(n4684), .Z(n5200) );
  OR2 U3285 ( .A(U7_DATA1_53), .B(n4662), .Z(n5199) );
  IV U3286 ( .A(n5201), .Z(n5197) );
  AN2 U3287 ( .A(n5202), .B(n5201), .Z(n5195) );
  OR2 U3288 ( .A(n5203), .B(n5204), .Z(n5201) );
  OR2 U3289 ( .A(n279), .B(n5205), .Z(n5204) );
  AN2 U3290 ( .A(ENCODER_DATA_IN[34]), .B(n4445), .Z(n5205) );
  AN2 U3291 ( .A(U24_Z_0), .B(n4446), .Z(n5203) );
  OR2 U3292 ( .A(n5206), .B(n5207), .Z(n5202) );
  AN2 U3293 ( .A(U7_DATA1_34), .B(n4684), .Z(n5207) );
  IV U3294 ( .A(U7_DATA1_53), .Z(n4684) );
  AN2 U3295 ( .A(U7_DATA1_53), .B(n4662), .Z(n5206) );
  IV U3296 ( .A(U7_DATA1_34), .Z(n4662) );
  AN2 U3297 ( .A(TEST_PAT_SEED_A[28]), .B(n4391), .Z(n5192) );
  AN2 U3298 ( .A(TEST_PAT_SEED_B[28]), .B(n4392), .Z(n5190) );
  OR2 U3299 ( .A(n5208), .B(n5209), .Z(U5_Z_27) );
  OR2 U3300 ( .A(n5210), .B(n5211), .Z(n5209) );
  OR2 U3301 ( .A(n5212), .B(n5213), .Z(n5211) );
  AN2 U3302 ( .A(U7_DATA4_27), .B(n4384), .Z(n5213) );
  AN2 U3303 ( .A(U7_DATA6_27), .B(n4385), .Z(n5212) );
  AN2 U3304 ( .A(n2661), .B(U7_DATA1_27), .Z(n5210) );
  OR2 U3305 ( .A(n5214), .B(n5215), .Z(n5208) );
  OR2 U3306 ( .A(n5216), .B(n5217), .Z(n5215) );
  AN2 U3307 ( .A(ENCODER_DATA_OUT[35]), .B(n4390), .Z(n5217) );
  IV U3308 ( .A(n5218), .Z(ENCODER_DATA_OUT[35]) );
  OR2 U3309 ( .A(n5219), .B(n5220), .Z(n5218) );
  AN2 U3310 ( .A(n5221), .B(n5222), .Z(n5220) );
  AN2 U3311 ( .A(n5223), .B(n5224), .Z(n5222) );
  OR2 U3312 ( .A(U7_DATA1_33), .B(n4718), .Z(n5224) );
  OR2 U3313 ( .A(U7_DATA1_52), .B(n4696), .Z(n5223) );
  IV U3314 ( .A(n5225), .Z(n5221) );
  AN2 U3315 ( .A(n5226), .B(n5225), .Z(n5219) );
  OR2 U3316 ( .A(n5227), .B(n5228), .Z(n5225) );
  OR2 U3317 ( .A(n279), .B(n5229), .Z(n5228) );
  AN2 U3318 ( .A(ENCODER_DATA_IN[33]), .B(n4445), .Z(n5229) );
  AN2 U3319 ( .A(U25_Z_1), .B(n4446), .Z(n5227) );
  OR2 U3320 ( .A(n5230), .B(n5231), .Z(n5226) );
  AN2 U3321 ( .A(U7_DATA1_33), .B(n4718), .Z(n5231) );
  IV U3322 ( .A(U7_DATA1_52), .Z(n4718) );
  AN2 U3323 ( .A(U7_DATA1_52), .B(n4696), .Z(n5230) );
  IV U3324 ( .A(U7_DATA1_33), .Z(n4696) );
  AN2 U3325 ( .A(TEST_PAT_SEED_A[27]), .B(n4391), .Z(n5216) );
  AN2 U3326 ( .A(TEST_PAT_SEED_B[27]), .B(n4392), .Z(n5214) );
  OR2 U3327 ( .A(n5232), .B(n5233), .Z(U5_Z_26) );
  OR2 U3328 ( .A(n5234), .B(n5235), .Z(n5233) );
  OR2 U3329 ( .A(n5236), .B(n5237), .Z(n5235) );
  AN2 U3330 ( .A(U7_DATA4_26), .B(n4384), .Z(n5237) );
  AN2 U3331 ( .A(U7_DATA6_26), .B(n4385), .Z(n5236) );
  AN2 U3332 ( .A(n2661), .B(U7_DATA1_26), .Z(n5234) );
  OR2 U3333 ( .A(n5238), .B(n5239), .Z(n5232) );
  OR2 U3334 ( .A(n5240), .B(n5241), .Z(n5239) );
  AN2 U3335 ( .A(ENCODER_DATA_OUT[34]), .B(n4390), .Z(n5241) );
  IV U3336 ( .A(n5242), .Z(ENCODER_DATA_OUT[34]) );
  OR2 U3337 ( .A(n5243), .B(n5244), .Z(n5242) );
  AN2 U3338 ( .A(n5245), .B(n5246), .Z(n5244) );
  AN2 U3339 ( .A(n5247), .B(n5248), .Z(n5246) );
  OR2 U3340 ( .A(U7_DATA1_32), .B(n4752), .Z(n5248) );
  OR2 U3341 ( .A(U7_DATA1_51), .B(n4730), .Z(n5247) );
  IV U3342 ( .A(n5249), .Z(n5245) );
  AN2 U3343 ( .A(n5250), .B(n5249), .Z(n5243) );
  OR2 U3344 ( .A(n5251), .B(n5252), .Z(n5249) );
  OR2 U3345 ( .A(n279), .B(n5253), .Z(n5252) );
  AN2 U3346 ( .A(ENCODER_DATA_IN[32]), .B(n4445), .Z(n5253) );
  AN2 U3347 ( .A(U25_Z_0), .B(n4446), .Z(n5251) );
  OR2 U3348 ( .A(n5254), .B(n5255), .Z(n5250) );
  AN2 U3349 ( .A(U7_DATA1_32), .B(n4752), .Z(n5255) );
  IV U3350 ( .A(U7_DATA1_51), .Z(n4752) );
  AN2 U3351 ( .A(U7_DATA1_51), .B(n4730), .Z(n5254) );
  IV U3352 ( .A(U7_DATA1_32), .Z(n4730) );
  AN2 U3353 ( .A(TEST_PAT_SEED_A[26]), .B(n4391), .Z(n5240) );
  AN2 U3354 ( .A(TEST_PAT_SEED_B[26]), .B(n4392), .Z(n5238) );
  OR2 U3355 ( .A(n5256), .B(n5257), .Z(U5_Z_25) );
  OR2 U3356 ( .A(n5258), .B(n5259), .Z(n5257) );
  OR2 U3357 ( .A(n5260), .B(n5261), .Z(n5259) );
  AN2 U3358 ( .A(U7_DATA4_25), .B(n4384), .Z(n5261) );
  AN2 U3359 ( .A(U7_DATA6_25), .B(n4385), .Z(n5260) );
  AN2 U3360 ( .A(n2661), .B(U7_DATA1_25), .Z(n5258) );
  OR2 U3361 ( .A(n5262), .B(n5263), .Z(n5256) );
  OR2 U3362 ( .A(n5264), .B(n5265), .Z(n5263) );
  AN2 U3363 ( .A(ENCODER_DATA_OUT[33]), .B(n4390), .Z(n5265) );
  IV U3364 ( .A(n5266), .Z(ENCODER_DATA_OUT[33]) );
  OR2 U3365 ( .A(n5267), .B(n5268), .Z(n5266) );
  AN2 U3366 ( .A(n5269), .B(n5270), .Z(n5268) );
  AN2 U3367 ( .A(n5271), .B(n5272), .Z(n5270) );
  OR2 U3368 ( .A(U7_DATA1_31), .B(n4786), .Z(n5272) );
  OR2 U3369 ( .A(U7_DATA1_50), .B(n4764), .Z(n5271) );
  IV U3370 ( .A(n5273), .Z(n5269) );
  AN2 U3371 ( .A(n5274), .B(n5273), .Z(n5267) );
  OR2 U3372 ( .A(n5275), .B(n5276), .Z(n5273) );
  OR2 U3373 ( .A(n279), .B(n5277), .Z(n5276) );
  AN2 U3374 ( .A(ENCODER_DATA_IN[31]), .B(n4445), .Z(n5277) );
  AN2 U3375 ( .A(U26_Z_2), .B(n4446), .Z(n5275) );
  OR2 U3376 ( .A(n5278), .B(n5279), .Z(n5274) );
  AN2 U3377 ( .A(U7_DATA1_31), .B(n4786), .Z(n5279) );
  IV U3378 ( .A(U7_DATA1_50), .Z(n4786) );
  AN2 U3379 ( .A(U7_DATA1_50), .B(n4764), .Z(n5278) );
  IV U3380 ( .A(U7_DATA1_31), .Z(n4764) );
  AN2 U3381 ( .A(TEST_PAT_SEED_A[25]), .B(n4391), .Z(n5264) );
  AN2 U3382 ( .A(TEST_PAT_SEED_B[25]), .B(n4392), .Z(n5262) );
  OR2 U3383 ( .A(n5280), .B(n5281), .Z(U5_Z_24) );
  OR2 U3384 ( .A(n5282), .B(n5283), .Z(n5281) );
  OR2 U3385 ( .A(n5284), .B(n5285), .Z(n5283) );
  AN2 U3386 ( .A(U7_DATA4_24), .B(n4384), .Z(n5285) );
  AN2 U3387 ( .A(U7_DATA6_24), .B(n4385), .Z(n5284) );
  AN2 U3388 ( .A(n2661), .B(U7_DATA1_24), .Z(n5282) );
  OR2 U3389 ( .A(n5286), .B(n5287), .Z(n5280) );
  OR2 U3390 ( .A(n5288), .B(n5289), .Z(n5287) );
  AN2 U3391 ( .A(ENCODER_DATA_OUT[32]), .B(n4390), .Z(n5289) );
  IV U3392 ( .A(n5290), .Z(ENCODER_DATA_OUT[32]) );
  OR2 U3393 ( .A(n5291), .B(n5292), .Z(n5290) );
  AN2 U3394 ( .A(n5293), .B(n5294), .Z(n5292) );
  AN2 U3395 ( .A(n5295), .B(n5296), .Z(n5294) );
  OR2 U3396 ( .A(U7_DATA1_30), .B(n4820), .Z(n5296) );
  OR2 U3397 ( .A(U7_DATA1_49), .B(n4798), .Z(n5295) );
  IV U3398 ( .A(n5297), .Z(n5293) );
  AN2 U3399 ( .A(n5298), .B(n5297), .Z(n5291) );
  OR2 U3400 ( .A(n5299), .B(n5300), .Z(n5297) );
  OR2 U3401 ( .A(n279), .B(n5301), .Z(n5300) );
  AN2 U3402 ( .A(ENCODER_DATA_IN[30]), .B(n4445), .Z(n5301) );
  AN2 U3403 ( .A(U26_Z_1), .B(n4446), .Z(n5299) );
  OR2 U3404 ( .A(n5302), .B(n5303), .Z(n5298) );
  AN2 U3405 ( .A(U7_DATA1_30), .B(n4820), .Z(n5303) );
  IV U3406 ( .A(U7_DATA1_49), .Z(n4820) );
  AN2 U3407 ( .A(U7_DATA1_49), .B(n4798), .Z(n5302) );
  IV U3408 ( .A(U7_DATA1_30), .Z(n4798) );
  AN2 U3409 ( .A(TEST_PAT_SEED_A[24]), .B(n4391), .Z(n5288) );
  AN2 U3410 ( .A(TEST_PAT_SEED_B[24]), .B(n4392), .Z(n5286) );
  OR2 U3411 ( .A(n5304), .B(n5305), .Z(U5_Z_23) );
  OR2 U3412 ( .A(n5306), .B(n5307), .Z(n5305) );
  OR2 U3413 ( .A(n5308), .B(n5309), .Z(n5307) );
  AN2 U3414 ( .A(U7_DATA4_23), .B(n4384), .Z(n5309) );
  AN2 U3415 ( .A(U7_DATA6_23), .B(n4385), .Z(n5308) );
  AN2 U3416 ( .A(n2661), .B(U7_DATA1_23), .Z(n5306) );
  OR2 U3417 ( .A(n5310), .B(n5311), .Z(n5304) );
  OR2 U3418 ( .A(n5312), .B(n5313), .Z(n5311) );
  AN2 U3419 ( .A(ENCODER_DATA_OUT[31]), .B(n4390), .Z(n5313) );
  IV U3420 ( .A(n5314), .Z(ENCODER_DATA_OUT[31]) );
  OR2 U3421 ( .A(n5315), .B(n5316), .Z(n5314) );
  AN2 U3422 ( .A(n5317), .B(n5318), .Z(n5316) );
  AN2 U3423 ( .A(n5319), .B(n5320), .Z(n5318) );
  OR2 U3424 ( .A(U7_DATA1_29), .B(n4842), .Z(n5320) );
  OR2 U3425 ( .A(U7_DATA1_48), .B(n4908), .Z(n5319) );
  IV U3426 ( .A(n5321), .Z(n5317) );
  AN2 U3427 ( .A(n5322), .B(n5321), .Z(n5315) );
  OR2 U3428 ( .A(n5323), .B(n5324), .Z(n5321) );
  OR2 U3429 ( .A(n279), .B(n5325), .Z(n5324) );
  AN2 U3430 ( .A(ENCODER_DATA_IN[29]), .B(n4445), .Z(n5325) );
  AN2 U3431 ( .A(U26_Z_0), .B(n4446), .Z(n5323) );
  OR2 U3432 ( .A(n5326), .B(n5327), .Z(n5322) );
  AN2 U3433 ( .A(U7_DATA1_29), .B(n4842), .Z(n5327) );
  IV U3434 ( .A(U7_DATA1_48), .Z(n4842) );
  AN2 U3435 ( .A(U7_DATA1_48), .B(n4908), .Z(n5326) );
  IV U3436 ( .A(U7_DATA1_29), .Z(n4908) );
  AN2 U3437 ( .A(TEST_PAT_SEED_A[23]), .B(n4391), .Z(n5312) );
  AN2 U3438 ( .A(TEST_PAT_SEED_B[23]), .B(n4392), .Z(n5310) );
  OR2 U3439 ( .A(n5328), .B(n5329), .Z(U5_Z_22) );
  OR2 U3440 ( .A(n5330), .B(n5331), .Z(n5329) );
  OR2 U3441 ( .A(n5332), .B(n5333), .Z(n5331) );
  AN2 U3442 ( .A(U7_DATA4_22), .B(n4384), .Z(n5333) );
  AN2 U3443 ( .A(U7_DATA6_22), .B(n4385), .Z(n5332) );
  AN2 U3444 ( .A(n2661), .B(U7_DATA1_22), .Z(n5330) );
  OR2 U3445 ( .A(n5334), .B(n5335), .Z(n5328) );
  OR2 U3446 ( .A(n5336), .B(n5337), .Z(n5335) );
  AN2 U3447 ( .A(ENCODER_DATA_OUT[30]), .B(n4390), .Z(n5337) );
  IV U3448 ( .A(n5338), .Z(ENCODER_DATA_OUT[30]) );
  OR2 U3449 ( .A(n5339), .B(n5340), .Z(n5338) );
  AN2 U3450 ( .A(n5341), .B(n5342), .Z(n5340) );
  AN2 U3451 ( .A(n5343), .B(n5344), .Z(n5342) );
  OR2 U3452 ( .A(U7_DATA1_28), .B(n4864), .Z(n5344) );
  OR2 U3453 ( .A(U7_DATA1_47), .B(n5155), .Z(n5343) );
  IV U3454 ( .A(n5345), .Z(n5341) );
  AN2 U3455 ( .A(n5346), .B(n5345), .Z(n5339) );
  OR2 U3456 ( .A(n5347), .B(n5348), .Z(n5345) );
  OR2 U3457 ( .A(n279), .B(n5349), .Z(n5348) );
  AN2 U3458 ( .A(ENCODER_DATA_IN[28]), .B(n4445), .Z(n5349) );
  AN2 U3459 ( .A(U27_Z_1), .B(n4446), .Z(n5347) );
  OR2 U3460 ( .A(n5350), .B(n5351), .Z(n5346) );
  AN2 U3461 ( .A(U7_DATA1_28), .B(n4864), .Z(n5351) );
  IV U3462 ( .A(U7_DATA1_47), .Z(n4864) );
  AN2 U3463 ( .A(U7_DATA1_47), .B(n5155), .Z(n5350) );
  IV U3464 ( .A(U7_DATA1_28), .Z(n5155) );
  AN2 U3465 ( .A(TEST_PAT_SEED_A[22]), .B(n4391), .Z(n5336) );
  AN2 U3466 ( .A(TEST_PAT_SEED_B[22]), .B(n4392), .Z(n5334) );
  OR2 U3467 ( .A(n5352), .B(n5353), .Z(U5_Z_21) );
  OR2 U3468 ( .A(n5354), .B(n5355), .Z(n5353) );
  OR2 U3469 ( .A(n5356), .B(n5357), .Z(n5355) );
  AN2 U3470 ( .A(U7_DATA4_21), .B(n4384), .Z(n5357) );
  AN2 U3471 ( .A(U7_DATA6_21), .B(n4385), .Z(n5356) );
  AN2 U3472 ( .A(n2661), .B(U7_DATA1_21), .Z(n5354) );
  OR2 U3473 ( .A(n5358), .B(n5359), .Z(n5352) );
  OR2 U3474 ( .A(n5360), .B(n5361), .Z(n5359) );
  AN2 U3475 ( .A(ENCODER_DATA_OUT[29]), .B(n4390), .Z(n5361) );
  IV U3476 ( .A(n5362), .Z(ENCODER_DATA_OUT[29]) );
  OR2 U3477 ( .A(n5363), .B(n5364), .Z(n5362) );
  AN2 U3478 ( .A(n5365), .B(n5366), .Z(n5364) );
  AN2 U3479 ( .A(n5367), .B(n5368), .Z(n5366) );
  OR2 U3480 ( .A(U7_DATA1_27), .B(n4886), .Z(n5368) );
  OR2 U3481 ( .A(U7_DATA1_46), .B(n5369), .Z(n5367) );
  IV U3482 ( .A(n5370), .Z(n5365) );
  AN2 U3483 ( .A(n5371), .B(n5370), .Z(n5363) );
  OR2 U3484 ( .A(n5372), .B(n5373), .Z(n5370) );
  OR2 U3485 ( .A(n279), .B(n5374), .Z(n5373) );
  AN2 U3486 ( .A(ENCODER_DATA_IN[27]), .B(n4445), .Z(n5374) );
  AN2 U3487 ( .A(U27_Z_0), .B(n4446), .Z(n5372) );
  OR2 U3488 ( .A(n5375), .B(n5376), .Z(n5371) );
  AN2 U3489 ( .A(U7_DATA1_27), .B(n4886), .Z(n5376) );
  IV U3490 ( .A(U7_DATA1_46), .Z(n4886) );
  AN2 U3491 ( .A(U7_DATA1_46), .B(n5369), .Z(n5375) );
  AN2 U3492 ( .A(TEST_PAT_SEED_A[21]), .B(n4391), .Z(n5360) );
  AN2 U3493 ( .A(TEST_PAT_SEED_B[21]), .B(n4392), .Z(n5358) );
  OR2 U3494 ( .A(n5377), .B(n5378), .Z(U5_Z_20) );
  OR2 U3495 ( .A(n5379), .B(n5380), .Z(n5378) );
  OR2 U3496 ( .A(n5381), .B(n5382), .Z(n5380) );
  AN2 U3497 ( .A(U7_DATA4_20), .B(n4384), .Z(n5382) );
  AN2 U3498 ( .A(U7_DATA6_20), .B(n4385), .Z(n5381) );
  AN2 U3499 ( .A(n2661), .B(U7_DATA1_20), .Z(n5379) );
  OR2 U3500 ( .A(n5383), .B(n5384), .Z(n5377) );
  OR2 U3501 ( .A(n5385), .B(n5386), .Z(n5384) );
  AN2 U3502 ( .A(ENCODER_DATA_OUT[28]), .B(n4390), .Z(n5386) );
  IV U3503 ( .A(n5387), .Z(ENCODER_DATA_OUT[28]) );
  OR2 U3504 ( .A(n5388), .B(n5389), .Z(n5387) );
  AN2 U3505 ( .A(n5390), .B(n5391), .Z(n5389) );
  AN2 U3506 ( .A(n5392), .B(n5393), .Z(n5391) );
  OR2 U3507 ( .A(U7_DATA1_26), .B(n4930), .Z(n5393) );
  OR2 U3508 ( .A(U7_DATA1_45), .B(n5394), .Z(n5392) );
  IV U3509 ( .A(n5395), .Z(n5390) );
  AN2 U3510 ( .A(n5396), .B(n5395), .Z(n5388) );
  OR2 U3511 ( .A(n5397), .B(n5398), .Z(n5395) );
  OR2 U3512 ( .A(n279), .B(n5399), .Z(n5398) );
  AN2 U3513 ( .A(ENCODER_DATA_IN[26]), .B(n4445), .Z(n5399) );
  AN2 U3514 ( .A(U28_Z_2), .B(n4446), .Z(n5397) );
  OR2 U3515 ( .A(n5400), .B(n5401), .Z(n5396) );
  AN2 U3516 ( .A(U7_DATA1_26), .B(n4930), .Z(n5401) );
  IV U3517 ( .A(U7_DATA1_45), .Z(n4930) );
  AN2 U3518 ( .A(U7_DATA1_45), .B(n5394), .Z(n5400) );
  AN2 U3519 ( .A(TEST_PAT_SEED_A[20]), .B(n4391), .Z(n5385) );
  AN2 U3520 ( .A(TEST_PAT_SEED_B[20]), .B(n4392), .Z(n5383) );
  OR2 U3521 ( .A(n5402), .B(n5403), .Z(U5_Z_2) );
  OR2 U3522 ( .A(n5404), .B(n5405), .Z(n5403) );
  OR2 U3523 ( .A(n5406), .B(n5407), .Z(n5405) );
  AN2 U3524 ( .A(U7_DATA4_2), .B(n4384), .Z(n5407) );
  AN2 U3525 ( .A(U7_DATA6_2), .B(n4385), .Z(n5406) );
  AN2 U3526 ( .A(n2661), .B(U7_DATA1_2), .Z(n5404) );
  OR2 U3527 ( .A(n5408), .B(n5409), .Z(n5402) );
  OR2 U3528 ( .A(n5410), .B(n5411), .Z(n5409) );
  AN2 U3529 ( .A(n4390), .B(ENCODER_DATA_OUT[10]), .Z(n5411) );
  AN2 U3530 ( .A(n5412), .B(n5413), .Z(ENCODER_DATA_OUT[10]) );
  IV U3531 ( .A(n5414), .Z(n5413) );
  AN2 U3532 ( .A(n5415), .B(n5416), .Z(n5414) );
  OR2 U3533 ( .A(n5416), .B(n5415), .Z(n5412) );
  OR2 U3534 ( .A(n5417), .B(n5418), .Z(n5415) );
  AN2 U3535 ( .A(U7_DATA1_27), .B(n5419), .Z(n5418) );
  IV U3536 ( .A(U7_DATA1_8), .Z(n5419) );
  AN2 U3537 ( .A(U7_DATA1_8), .B(n5369), .Z(n5417) );
  IV U3538 ( .A(U7_DATA1_27), .Z(n5369) );
  OR2 U3539 ( .A(n5420), .B(n5421), .Z(n5416) );
  OR2 U3540 ( .A(n279), .B(n5422), .Z(n5421) );
  AN2 U3541 ( .A(ENCODER_DATA_IN[8]), .B(n4445), .Z(n5422) );
  AN2 U3542 ( .A(U34_Z_0), .B(n4446), .Z(n5420) );
  AN2 U3543 ( .A(TEST_PAT_SEED_A[2]), .B(n4391), .Z(n5410) );
  AN2 U3544 ( .A(TEST_PAT_SEED_B[2]), .B(n4392), .Z(n5408) );
  OR2 U3545 ( .A(n5423), .B(n5424), .Z(U5_Z_19) );
  OR2 U3546 ( .A(n5425), .B(n5426), .Z(n5424) );
  OR2 U3547 ( .A(n5427), .B(n5428), .Z(n5426) );
  AN2 U3548 ( .A(U7_DATA4_19), .B(n4384), .Z(n5428) );
  AN2 U3549 ( .A(U7_DATA6_19), .B(n4385), .Z(n5427) );
  AN2 U3550 ( .A(n2661), .B(U7_DATA1_19), .Z(n5425) );
  OR2 U3551 ( .A(n5429), .B(n5430), .Z(n5423) );
  OR2 U3552 ( .A(n5431), .B(n5432), .Z(n5430) );
  AN2 U3553 ( .A(ENCODER_DATA_OUT[27]), .B(n4390), .Z(n5432) );
  IV U3554 ( .A(n5433), .Z(ENCODER_DATA_OUT[27]) );
  OR2 U3555 ( .A(n5434), .B(n5435), .Z(n5433) );
  AN2 U3556 ( .A(n5436), .B(n5437), .Z(n5435) );
  AN2 U3557 ( .A(n5438), .B(n5439), .Z(n5437) );
  OR2 U3558 ( .A(U7_DATA1_25), .B(n4952), .Z(n5439) );
  OR2 U3559 ( .A(U7_DATA1_44), .B(n5440), .Z(n5438) );
  IV U3560 ( .A(n5441), .Z(n5436) );
  AN2 U3561 ( .A(n5442), .B(n5441), .Z(n5434) );
  OR2 U3562 ( .A(n5443), .B(n5444), .Z(n5441) );
  OR2 U3563 ( .A(n279), .B(n5445), .Z(n5444) );
  AN2 U3564 ( .A(ENCODER_DATA_IN[25]), .B(n4445), .Z(n5445) );
  AN2 U3565 ( .A(U28_Z_1), .B(n4446), .Z(n5443) );
  OR2 U3566 ( .A(n5446), .B(n5447), .Z(n5442) );
  AN2 U3567 ( .A(U7_DATA1_25), .B(n4952), .Z(n5447) );
  IV U3568 ( .A(U7_DATA1_44), .Z(n4952) );
  AN2 U3569 ( .A(U7_DATA1_44), .B(n5440), .Z(n5446) );
  AN2 U3570 ( .A(TEST_PAT_SEED_A[19]), .B(n4391), .Z(n5431) );
  AN2 U3571 ( .A(TEST_PAT_SEED_B[19]), .B(n4392), .Z(n5429) );
  OR2 U3572 ( .A(n5448), .B(n5449), .Z(U5_Z_18) );
  OR2 U3573 ( .A(n5450), .B(n5451), .Z(n5449) );
  OR2 U3574 ( .A(n5452), .B(n5453), .Z(n5451) );
  AN2 U3575 ( .A(U7_DATA4_18), .B(n4384), .Z(n5453) );
  AN2 U3576 ( .A(U7_DATA6_18), .B(n4385), .Z(n5452) );
  AN2 U3577 ( .A(n2661), .B(U7_DATA1_18), .Z(n5450) );
  OR2 U3578 ( .A(n5454), .B(n5455), .Z(n5448) );
  OR2 U3579 ( .A(n5456), .B(n5457), .Z(n5455) );
  AN2 U3580 ( .A(n4390), .B(ENCODER_DATA_OUT[26]), .Z(n5457) );
  IV U3581 ( .A(n4439), .Z(ENCODER_DATA_OUT[26]) );
  OR2 U3582 ( .A(n5458), .B(n5459), .Z(n4439) );
  AN2 U3583 ( .A(n5460), .B(n5461), .Z(n5459) );
  IV U3584 ( .A(n5462), .Z(n5458) );
  OR2 U3585 ( .A(n5461), .B(n5460), .Z(n5462) );
  OR2 U3586 ( .A(n5463), .B(n5464), .Z(n5460) );
  IV U3587 ( .A(n5465), .Z(n5464) );
  OR2 U3588 ( .A(n5466), .B(U7_DATA1_43), .Z(n5465) );
  AN2 U3589 ( .A(U7_DATA1_43), .B(n5466), .Z(n5463) );
  OR2 U3590 ( .A(n5467), .B(n5468), .Z(n5461) );
  OR2 U3591 ( .A(n281), .B(n5469), .Z(n5468) );
  AN2 U3592 ( .A(ENCODER_DATA_IN[24]), .B(n4445), .Z(n5469) );
  AN2 U3593 ( .A(U28_Z_0), .B(n4446), .Z(n5467) );
  AN2 U3594 ( .A(TEST_PAT_SEED_A[18]), .B(n4391), .Z(n5456) );
  AN2 U3595 ( .A(TEST_PAT_SEED_B[18]), .B(n4392), .Z(n5454) );
  OR2 U3596 ( .A(n5470), .B(n5471), .Z(U5_Z_17) );
  OR2 U3597 ( .A(n5472), .B(n5473), .Z(n5471) );
  OR2 U3598 ( .A(n5474), .B(n5475), .Z(n5473) );
  AN2 U3599 ( .A(U7_DATA4_17), .B(n4384), .Z(n5475) );
  AN2 U3600 ( .A(U7_DATA6_17), .B(n4385), .Z(n5474) );
  AN2 U3601 ( .A(n2661), .B(U7_DATA1_17), .Z(n5472) );
  OR2 U3602 ( .A(n5476), .B(n5477), .Z(n5470) );
  OR2 U3603 ( .A(n5478), .B(n5479), .Z(n5477) );
  AN2 U3604 ( .A(n4390), .B(ENCODER_DATA_OUT[25]), .Z(n5479) );
  AN2 U3605 ( .A(n5480), .B(n5481), .Z(ENCODER_DATA_OUT[25]) );
  IV U3606 ( .A(n5482), .Z(n5481) );
  AN2 U3607 ( .A(n5483), .B(n5484), .Z(n5482) );
  OR2 U3608 ( .A(n5484), .B(n5483), .Z(n5480) );
  OR2 U3609 ( .A(n5485), .B(n5486), .Z(n5483) );
  IV U3610 ( .A(n5487), .Z(n5486) );
  OR2 U3611 ( .A(n5488), .B(U7_DATA1_42), .Z(n5487) );
  AN2 U3612 ( .A(U7_DATA1_42), .B(n5488), .Z(n5485) );
  OR2 U3613 ( .A(n5489), .B(n5490), .Z(n5484) );
  OR2 U3614 ( .A(n279), .B(n5491), .Z(n5490) );
  AN2 U3615 ( .A(ENCODER_DATA_IN[23]), .B(n4445), .Z(n5491) );
  AN2 U3616 ( .A(U29_Z_1), .B(n4446), .Z(n5489) );
  AN2 U3617 ( .A(TEST_PAT_SEED_A[17]), .B(n4391), .Z(n5478) );
  AN2 U3618 ( .A(TEST_PAT_SEED_B[17]), .B(n4392), .Z(n5476) );
  OR2 U3619 ( .A(n5492), .B(n5493), .Z(U5_Z_16) );
  OR2 U3620 ( .A(n5494), .B(n5495), .Z(n5493) );
  OR2 U3621 ( .A(n5496), .B(n5497), .Z(n5495) );
  AN2 U3622 ( .A(U7_DATA4_16), .B(n4384), .Z(n5497) );
  AN2 U3623 ( .A(U7_DATA6_16), .B(n4385), .Z(n5496) );
  AN2 U3624 ( .A(n2661), .B(U7_DATA1_16), .Z(n5494) );
  OR2 U3625 ( .A(n5498), .B(n5499), .Z(n5492) );
  OR2 U3626 ( .A(n5500), .B(n5501), .Z(n5499) );
  AN2 U3627 ( .A(n4390), .B(ENCODER_DATA_OUT[24]), .Z(n5501) );
  AN2 U3628 ( .A(n5502), .B(n5503), .Z(ENCODER_DATA_OUT[24]) );
  IV U3629 ( .A(n5504), .Z(n5503) );
  AN2 U3630 ( .A(n5505), .B(n5506), .Z(n5504) );
  OR2 U3631 ( .A(n5506), .B(n5505), .Z(n5502) );
  OR2 U3632 ( .A(n5507), .B(n5508), .Z(n5505) );
  IV U3633 ( .A(n5509), .Z(n5508) );
  OR2 U3634 ( .A(n5510), .B(U7_DATA1_41), .Z(n5509) );
  AN2 U3635 ( .A(U7_DATA1_41), .B(n5510), .Z(n5507) );
  OR2 U3636 ( .A(n5511), .B(n5512), .Z(n5506) );
  OR2 U3637 ( .A(n279), .B(n5513), .Z(n5512) );
  AN2 U3638 ( .A(ENCODER_DATA_IN[22]), .B(n4445), .Z(n5513) );
  AN2 U3639 ( .A(U29_Z_0), .B(n4446), .Z(n5511) );
  AN2 U3640 ( .A(TEST_PAT_SEED_A[16]), .B(n4391), .Z(n5500) );
  AN2 U3641 ( .A(TEST_PAT_SEED_B[16]), .B(n4392), .Z(n5498) );
  OR2 U3642 ( .A(n5514), .B(n5515), .Z(U5_Z_15) );
  OR2 U3643 ( .A(n5516), .B(n5517), .Z(n5515) );
  OR2 U3644 ( .A(n5518), .B(n5519), .Z(n5517) );
  AN2 U3645 ( .A(U7_DATA4_15), .B(n4384), .Z(n5519) );
  AN2 U3646 ( .A(U7_DATA6_15), .B(n4385), .Z(n5518) );
  AN2 U3647 ( .A(n2661), .B(U7_DATA1_15), .Z(n5516) );
  OR2 U3648 ( .A(n5520), .B(n5521), .Z(n5514) );
  OR2 U3649 ( .A(n5522), .B(n5523), .Z(n5521) );
  AN2 U3650 ( .A(n4390), .B(ENCODER_DATA_OUT[23]), .Z(n5523) );
  AN2 U3651 ( .A(n5524), .B(n5525), .Z(ENCODER_DATA_OUT[23]) );
  IV U3652 ( .A(n5526), .Z(n5525) );
  AN2 U3653 ( .A(n5527), .B(n5528), .Z(n5526) );
  OR2 U3654 ( .A(n5528), .B(n5527), .Z(n5524) );
  OR2 U3655 ( .A(n5529), .B(n5530), .Z(n5527) );
  IV U3656 ( .A(n5531), .Z(n5530) );
  OR2 U3657 ( .A(n5532), .B(U7_DATA1_40), .Z(n5531) );
  AN2 U3658 ( .A(U7_DATA1_40), .B(n5532), .Z(n5529) );
  OR2 U3659 ( .A(n5533), .B(n5534), .Z(n5528) );
  OR2 U3660 ( .A(n279), .B(n5535), .Z(n5534) );
  AN2 U3661 ( .A(ENCODER_DATA_IN[21]), .B(n4445), .Z(n5535) );
  AN2 U3662 ( .A(U30_Z_1), .B(n4446), .Z(n5533) );
  AN2 U3663 ( .A(TEST_PAT_SEED_A[15]), .B(n4391), .Z(n5522) );
  AN2 U3664 ( .A(TEST_PAT_SEED_B[15]), .B(n4392), .Z(n5520) );
  OR2 U3665 ( .A(n5536), .B(n5537), .Z(U5_Z_14) );
  OR2 U3666 ( .A(n5538), .B(n5539), .Z(n5537) );
  OR2 U3667 ( .A(n5540), .B(n5541), .Z(n5539) );
  AN2 U3668 ( .A(U7_DATA4_14), .B(n4384), .Z(n5541) );
  AN2 U3669 ( .A(U7_DATA6_14), .B(n4385), .Z(n5540) );
  AN2 U3670 ( .A(n2661), .B(U7_DATA1_14), .Z(n5538) );
  OR2 U3671 ( .A(n5542), .B(n5543), .Z(n5536) );
  OR2 U3672 ( .A(n5544), .B(n5545), .Z(n5543) );
  AN2 U3673 ( .A(n4390), .B(ENCODER_DATA_OUT[22]), .Z(n5545) );
  AN2 U3674 ( .A(n5546), .B(n5547), .Z(ENCODER_DATA_OUT[22]) );
  IV U3675 ( .A(n5548), .Z(n5547) );
  AN2 U3676 ( .A(n5549), .B(n5550), .Z(n5548) );
  OR2 U3677 ( .A(n5550), .B(n5549), .Z(n5546) );
  OR2 U3678 ( .A(n5551), .B(n5552), .Z(n5549) );
  IV U3679 ( .A(n5553), .Z(n5552) );
  OR2 U3680 ( .A(n5554), .B(U7_DATA1_39), .Z(n5553) );
  AN2 U3681 ( .A(U7_DATA1_39), .B(n5554), .Z(n5551) );
  OR2 U3682 ( .A(n5555), .B(n5556), .Z(n5550) );
  OR2 U3683 ( .A(n279), .B(n5557), .Z(n5556) );
  AN2 U3684 ( .A(ENCODER_DATA_IN[20]), .B(n4445), .Z(n5557) );
  AN2 U3685 ( .A(U30_Z_0), .B(n4446), .Z(n5555) );
  AN2 U3686 ( .A(TEST_PAT_SEED_A[14]), .B(n4391), .Z(n5544) );
  AN2 U3687 ( .A(TEST_PAT_SEED_B[14]), .B(n4392), .Z(n5542) );
  OR2 U3688 ( .A(n5558), .B(n5559), .Z(U5_Z_13) );
  OR2 U3689 ( .A(n5560), .B(n5561), .Z(n5559) );
  OR2 U3690 ( .A(n5562), .B(n5563), .Z(n5561) );
  AN2 U3691 ( .A(U7_DATA4_13), .B(n4384), .Z(n5563) );
  AN2 U3692 ( .A(U7_DATA6_13), .B(n4385), .Z(n5562) );
  AN2 U3693 ( .A(n2661), .B(U7_DATA1_13), .Z(n5560) );
  OR2 U3694 ( .A(n5564), .B(n5565), .Z(n5558) );
  OR2 U3695 ( .A(n5566), .B(n5567), .Z(n5565) );
  AN2 U3696 ( .A(n4390), .B(ENCODER_DATA_OUT[21]), .Z(n5567) );
  AN2 U3697 ( .A(n5568), .B(n5569), .Z(ENCODER_DATA_OUT[21]) );
  IV U3698 ( .A(n5570), .Z(n5569) );
  AN2 U3699 ( .A(n5571), .B(n5572), .Z(n5570) );
  OR2 U3700 ( .A(n5572), .B(n5571), .Z(n5568) );
  OR2 U3701 ( .A(n5573), .B(n5574), .Z(n5571) );
  AN2 U3702 ( .A(U7_DATA1_19), .B(n5079), .Z(n5574) );
  IV U3703 ( .A(U7_DATA1_38), .Z(n5079) );
  AN2 U3704 ( .A(U7_DATA1_38), .B(n5575), .Z(n5573) );
  OR2 U3705 ( .A(n5576), .B(n5577), .Z(n5572) );
  OR2 U3706 ( .A(n279), .B(n5578), .Z(n5577) );
  AN2 U3707 ( .A(ENCODER_DATA_IN[19]), .B(n4445), .Z(n5578) );
  AN2 U3708 ( .A(U31_Z_3), .B(n4446), .Z(n5576) );
  AN2 U3709 ( .A(TEST_PAT_SEED_A[13]), .B(n4391), .Z(n5566) );
  AN2 U3710 ( .A(TEST_PAT_SEED_B[13]), .B(n4392), .Z(n5564) );
  OR2 U3711 ( .A(n5579), .B(n5580), .Z(U5_Z_12) );
  OR2 U3712 ( .A(n5581), .B(n5582), .Z(n5580) );
  OR2 U3713 ( .A(n5583), .B(n5584), .Z(n5582) );
  AN2 U3714 ( .A(U7_DATA4_12), .B(n4384), .Z(n5584) );
  AN2 U3715 ( .A(U7_DATA6_12), .B(n4385), .Z(n5583) );
  AN2 U3716 ( .A(n2661), .B(U7_DATA1_12), .Z(n5581) );
  OR2 U3717 ( .A(n5585), .B(n5586), .Z(n5579) );
  OR2 U3718 ( .A(n5587), .B(n5588), .Z(n5586) );
  AN2 U3719 ( .A(n4390), .B(ENCODER_DATA_OUT[20]), .Z(n5588) );
  AN2 U3720 ( .A(n5589), .B(n5590), .Z(ENCODER_DATA_OUT[20]) );
  IV U3721 ( .A(n5591), .Z(n5590) );
  AN2 U3722 ( .A(n5592), .B(n5593), .Z(n5591) );
  OR2 U3723 ( .A(n5593), .B(n5592), .Z(n5589) );
  OR2 U3724 ( .A(n5594), .B(n5595), .Z(n5592) );
  AN2 U3725 ( .A(U7_DATA1_18), .B(n5104), .Z(n5595) );
  IV U3726 ( .A(U7_DATA1_37), .Z(n5104) );
  AN2 U3727 ( .A(U7_DATA1_37), .B(n5596), .Z(n5594) );
  IV U3728 ( .A(U7_DATA1_18), .Z(n5596) );
  OR2 U3729 ( .A(n5597), .B(n5598), .Z(n5593) );
  OR2 U3730 ( .A(n279), .B(n5599), .Z(n5598) );
  AN2 U3731 ( .A(ENCODER_DATA_IN[18]), .B(n4445), .Z(n5599) );
  AN2 U3732 ( .A(U31_Z_2), .B(n4446), .Z(n5597) );
  AN2 U3733 ( .A(TEST_PAT_SEED_A[12]), .B(n4391), .Z(n5587) );
  AN2 U3734 ( .A(TEST_PAT_SEED_B[12]), .B(n4392), .Z(n5585) );
  OR2 U3735 ( .A(n5600), .B(n5601), .Z(U5_Z_11) );
  OR2 U3736 ( .A(n5602), .B(n5603), .Z(n5601) );
  OR2 U3737 ( .A(n5604), .B(n5605), .Z(n5603) );
  AN2 U3738 ( .A(U7_DATA4_11), .B(n4384), .Z(n5605) );
  AN2 U3739 ( .A(U7_DATA6_11), .B(n4385), .Z(n5604) );
  AN2 U3740 ( .A(n2661), .B(U7_DATA1_11), .Z(n5602) );
  OR2 U3741 ( .A(n5606), .B(n5607), .Z(n5600) );
  OR2 U3742 ( .A(n5608), .B(n5609), .Z(n5607) );
  AN2 U3743 ( .A(n4390), .B(ENCODER_DATA_OUT[19]), .Z(n5609) );
  AN2 U3744 ( .A(n5610), .B(n5611), .Z(ENCODER_DATA_OUT[19]) );
  IV U3745 ( .A(n5612), .Z(n5611) );
  AN2 U3746 ( .A(n5613), .B(n5614), .Z(n5612) );
  OR2 U3747 ( .A(n5614), .B(n5613), .Z(n5610) );
  OR2 U3748 ( .A(n5615), .B(n5616), .Z(n5613) );
  AN2 U3749 ( .A(U7_DATA1_17), .B(n5129), .Z(n5616) );
  IV U3750 ( .A(U7_DATA1_36), .Z(n5129) );
  AN2 U3751 ( .A(U7_DATA1_36), .B(n5617), .Z(n5615) );
  IV U3752 ( .A(U7_DATA1_17), .Z(n5617) );
  OR2 U3753 ( .A(n5618), .B(n5619), .Z(n5614) );
  OR2 U3754 ( .A(n279), .B(n5620), .Z(n5619) );
  AN2 U3755 ( .A(ENCODER_DATA_IN[17]), .B(n4445), .Z(n5620) );
  AN2 U3756 ( .A(U31_Z_1), .B(n4446), .Z(n5618) );
  AN2 U3757 ( .A(TEST_PAT_SEED_A[11]), .B(n4391), .Z(n5608) );
  AN2 U3758 ( .A(TEST_PAT_SEED_B[11]), .B(n4392), .Z(n5606) );
  OR2 U3759 ( .A(n5621), .B(n5622), .Z(U5_Z_10) );
  OR2 U3760 ( .A(n5623), .B(n5624), .Z(n5622) );
  OR2 U3761 ( .A(n5625), .B(n5626), .Z(n5624) );
  AN2 U3762 ( .A(U7_DATA4_10), .B(n4384), .Z(n5626) );
  AN2 U3763 ( .A(U7_DATA6_10), .B(n4385), .Z(n5625) );
  AN2 U3764 ( .A(n2661), .B(U7_DATA1_10), .Z(n5623) );
  OR2 U3765 ( .A(n5627), .B(n5628), .Z(n5621) );
  OR2 U3766 ( .A(n5629), .B(n5630), .Z(n5628) );
  AN2 U3767 ( .A(n4390), .B(ENCODER_DATA_OUT[18]), .Z(n5630) );
  AN2 U3768 ( .A(n5631), .B(n5632), .Z(ENCODER_DATA_OUT[18]) );
  IV U3769 ( .A(n5633), .Z(n5632) );
  AN2 U3770 ( .A(n5634), .B(n5635), .Z(n5633) );
  OR2 U3771 ( .A(n5635), .B(n5634), .Z(n5631) );
  OR2 U3772 ( .A(n5636), .B(n5637), .Z(n5634) );
  AN2 U3773 ( .A(U7_DATA1_16), .B(n5176), .Z(n5637) );
  IV U3774 ( .A(U7_DATA1_35), .Z(n5176) );
  AN2 U3775 ( .A(U7_DATA1_35), .B(n5638), .Z(n5636) );
  IV U3776 ( .A(U7_DATA1_16), .Z(n5638) );
  OR2 U3777 ( .A(n5639), .B(n5640), .Z(n5635) );
  OR2 U3778 ( .A(n279), .B(n5641), .Z(n5640) );
  AN2 U3779 ( .A(ENCODER_DATA_IN[16]), .B(n4445), .Z(n5641) );
  AN2 U3780 ( .A(U31_Z_0), .B(n4446), .Z(n5639) );
  AN2 U3781 ( .A(TEST_PAT_SEED_A[10]), .B(n4391), .Z(n5629) );
  AN2 U3782 ( .A(TEST_PAT_SEED_B[10]), .B(n4392), .Z(n5627) );
  OR2 U3783 ( .A(n5642), .B(n5643), .Z(U5_Z_1) );
  OR2 U3784 ( .A(n5644), .B(n5645), .Z(n5643) );
  OR2 U3785 ( .A(n5646), .B(n5647), .Z(n5645) );
  AN2 U3786 ( .A(U7_DATA4_1), .B(n4384), .Z(n5647) );
  AN2 U3787 ( .A(U7_DATA6_1), .B(n4385), .Z(n5646) );
  AN2 U3788 ( .A(n2661), .B(U7_DATA1_1), .Z(n5644) );
  OR2 U3789 ( .A(n5648), .B(n5649), .Z(n5642) );
  OR2 U3790 ( .A(n5650), .B(n5651), .Z(n5649) );
  AN2 U3791 ( .A(n4390), .B(ENCODER_DATA_OUT[9]), .Z(n5651) );
  AN2 U3792 ( .A(n5652), .B(n5653), .Z(ENCODER_DATA_OUT[9]) );
  IV U3793 ( .A(n5654), .Z(n5653) );
  AN2 U3794 ( .A(n5655), .B(n5656), .Z(n5654) );
  OR2 U3795 ( .A(n5656), .B(n5655), .Z(n5652) );
  OR2 U3796 ( .A(n5657), .B(n5658), .Z(n5655) );
  AN2 U3797 ( .A(U7_DATA1_26), .B(n5659), .Z(n5658) );
  IV U3798 ( .A(U7_DATA1_7), .Z(n5659) );
  AN2 U3799 ( .A(U7_DATA1_7), .B(n5394), .Z(n5657) );
  IV U3800 ( .A(U7_DATA1_26), .Z(n5394) );
  OR2 U3801 ( .A(n5660), .B(n5661), .Z(n5656) );
  OR2 U3802 ( .A(n279), .B(n5662), .Z(n5661) );
  AN2 U3803 ( .A(ENCODER_DATA_IN[7]), .B(n4445), .Z(n5662) );
  AN2 U3804 ( .A(U10_DATA2_7), .B(n4446), .Z(n5660) );
  AN2 U3805 ( .A(TEST_PAT_SEED_A[1]), .B(n4391), .Z(n5650) );
  AN2 U3806 ( .A(TEST_PAT_SEED_B[1]), .B(n4392), .Z(n5648) );
  OR2 U3807 ( .A(n5663), .B(n5664), .Z(U5_Z_0) );
  OR2 U3808 ( .A(n5665), .B(n5666), .Z(n5664) );
  OR2 U3809 ( .A(n5667), .B(n5668), .Z(n5666) );
  AN2 U3810 ( .A(U7_DATA4_0), .B(n4384), .Z(n5668) );
  AN2 U3811 ( .A(n5669), .B(n5670), .Z(n4384) );
  AN2 U3812 ( .A(U7_DATA6_0), .B(n4385), .Z(n5667) );
  AN2 U3813 ( .A(n5671), .B(n5672), .Z(n4385) );
  AN2 U3814 ( .A(n940), .B(n5670), .Z(n5672) );
  IV U3815 ( .A(n5673), .Z(n5671) );
  OR2 U3816 ( .A(n949), .B(n5669), .Z(n5673) );
  AN2 U3817 ( .A(n2661), .B(U7_DATA1_0), .Z(n5665) );
  OR2 U3818 ( .A(n5674), .B(n5675), .Z(n5663) );
  OR2 U3819 ( .A(n5676), .B(n5677), .Z(n5675) );
  AN2 U3820 ( .A(n4390), .B(ENCODER_DATA_OUT[8]), .Z(n5677) );
  AN2 U3821 ( .A(n5678), .B(n5679), .Z(ENCODER_DATA_OUT[8]) );
  IV U3822 ( .A(n5680), .Z(n5679) );
  AN2 U3823 ( .A(n5681), .B(n5682), .Z(n5680) );
  OR2 U3824 ( .A(n5682), .B(n5681), .Z(n5678) );
  OR2 U3825 ( .A(n5683), .B(n5684), .Z(n5681) );
  AN2 U3826 ( .A(U7_DATA1_25), .B(n5685), .Z(n5684) );
  IV U3827 ( .A(U7_DATA1_6), .Z(n5685) );
  AN2 U3828 ( .A(U7_DATA1_6), .B(n5440), .Z(n5683) );
  IV U3829 ( .A(U7_DATA1_25), .Z(n5440) );
  OR2 U3830 ( .A(n5686), .B(n5687), .Z(n5682) );
  OR2 U3831 ( .A(n281), .B(n5688), .Z(n5687) );
  AN2 U3832 ( .A(ENCODER_DATA_IN[6]), .B(n4445), .Z(n5688) );
  AN2 U3833 ( .A(U10_DATA2_6), .B(n4446), .Z(n5686) );
  AN2 U3834 ( .A(n967), .B(n278), .Z(n4390) );
  AN2 U3835 ( .A(TEST_PAT_SEED_A[0]), .B(n4391), .Z(n5676) );
  AN2 U3836 ( .A(n1970), .B(n5689), .Z(n4391) );
  IV U3837 ( .A(n5690), .Z(n5689) );
  OR2 U3838 ( .A(n919), .B(n3749), .Z(n5690) );
  AN2 U3839 ( .A(TEST_PAT_SEED_B[0]), .B(n4392), .Z(n5674) );
  AN2 U3840 ( .A(n5670), .B(n5691), .Z(n4392) );
  IV U3841 ( .A(n5692), .Z(n5691) );
  OR2 U3842 ( .A(n940), .B(n5669), .Z(n5692) );
  IV U3843 ( .A(n931), .Z(n5669) );
  AN2 U3844 ( .A(n919), .B(n5693), .Z(n5670) );
  AN2 U3845 ( .A(n5694), .B(n1970), .Z(n5693) );
  IV U3846 ( .A(n3749), .Z(n5694) );
  AN2 U3847 ( .A(n5695), .B(n5696), .Z(ENCODER_DATA_OUT[7]) );
  IV U3848 ( .A(n5697), .Z(n5696) );
  AN2 U3849 ( .A(n5698), .B(n5699), .Z(n5697) );
  OR2 U3850 ( .A(n5699), .B(n5698), .Z(n5695) );
  OR2 U3851 ( .A(n5700), .B(n5701), .Z(n5698) );
  AN2 U3852 ( .A(U7_DATA1_24), .B(n5702), .Z(n5701) );
  IV U3853 ( .A(U7_DATA1_5), .Z(n5702) );
  AN2 U3854 ( .A(U7_DATA1_5), .B(n5466), .Z(n5700) );
  IV U3855 ( .A(U7_DATA1_24), .Z(n5466) );
  OR2 U3856 ( .A(n5703), .B(n5704), .Z(n5699) );
  OR2 U3857 ( .A(n279), .B(n5705), .Z(n5704) );
  AN2 U3858 ( .A(ENCODER_DATA_IN[5]), .B(n4445), .Z(n5705) );
  AN2 U3859 ( .A(U10_DATA2_5), .B(n4446), .Z(n5703) );
  AN2 U3860 ( .A(n5706), .B(n5707), .Z(ENCODER_DATA_OUT[6]) );
  IV U3861 ( .A(n5708), .Z(n5707) );
  AN2 U3862 ( .A(n5709), .B(n5710), .Z(n5708) );
  OR2 U3863 ( .A(n5710), .B(n5709), .Z(n5706) );
  OR2 U3864 ( .A(n5711), .B(n5712), .Z(n5709) );
  AN2 U3865 ( .A(U7_DATA1_23), .B(n5713), .Z(n5712) );
  IV U3866 ( .A(U7_DATA1_4), .Z(n5713) );
  AN2 U3867 ( .A(U7_DATA1_4), .B(n5488), .Z(n5711) );
  IV U3868 ( .A(U7_DATA1_23), .Z(n5488) );
  OR2 U3869 ( .A(n5714), .B(n5715), .Z(n5710) );
  OR2 U3870 ( .A(n281), .B(n5716), .Z(n5715) );
  AN2 U3871 ( .A(ENCODER_DATA_IN[4]), .B(n4445), .Z(n5716) );
  AN2 U3872 ( .A(U10_DATA2_4), .B(n4446), .Z(n5714) );
  AN2 U3873 ( .A(n5717), .B(n5718), .Z(ENCODER_DATA_OUT[5]) );
  IV U3874 ( .A(n5719), .Z(n5718) );
  AN2 U3875 ( .A(n5720), .B(n5721), .Z(n5719) );
  OR2 U3876 ( .A(n5721), .B(n5720), .Z(n5717) );
  OR2 U3877 ( .A(n5722), .B(n5723), .Z(n5720) );
  AN2 U3878 ( .A(U7_DATA1_22), .B(n5724), .Z(n5723) );
  IV U3879 ( .A(U7_DATA1_3), .Z(n5724) );
  AN2 U3880 ( .A(U7_DATA1_3), .B(n5510), .Z(n5722) );
  IV U3881 ( .A(U7_DATA1_22), .Z(n5510) );
  OR2 U3882 ( .A(n5725), .B(n5726), .Z(n5721) );
  OR2 U3883 ( .A(n279), .B(n5727), .Z(n5726) );
  AN2 U3884 ( .A(ENCODER_DATA_IN[3]), .B(n4445), .Z(n5727) );
  AN2 U3885 ( .A(U10_DATA2_3), .B(n4446), .Z(n5725) );
  AN2 U3886 ( .A(n5728), .B(n5729), .Z(ENCODER_DATA_OUT[4]) );
  IV U3887 ( .A(n5730), .Z(n5729) );
  AN2 U3888 ( .A(n5731), .B(n5732), .Z(n5730) );
  OR2 U3889 ( .A(n5732), .B(n5731), .Z(n5728) );
  OR2 U3890 ( .A(n5733), .B(n5734), .Z(n5731) );
  AN2 U3891 ( .A(U7_DATA1_2), .B(n5532), .Z(n5734) );
  IV U3892 ( .A(U7_DATA1_21), .Z(n5532) );
  AN2 U3893 ( .A(U7_DATA1_21), .B(n5735), .Z(n5733) );
  IV U3894 ( .A(U7_DATA1_2), .Z(n5735) );
  OR2 U3895 ( .A(n5736), .B(n5737), .Z(n5732) );
  OR2 U3896 ( .A(n281), .B(n5738), .Z(n5737) );
  AN2 U3897 ( .A(ENCODER_DATA_IN[2]), .B(n4445), .Z(n5738) );
  AN2 U3898 ( .A(U10_DATA2_2), .B(n4446), .Z(n5736) );
  AN2 U3899 ( .A(n5739), .B(n5740), .Z(ENCODER_DATA_OUT[3]) );
  IV U3900 ( .A(n5741), .Z(n5740) );
  AN2 U3901 ( .A(n5742), .B(n5743), .Z(n5741) );
  OR2 U3902 ( .A(n5743), .B(n5742), .Z(n5739) );
  OR2 U3903 ( .A(n5744), .B(n5745), .Z(n5742) );
  AN2 U3904 ( .A(U7_DATA1_1), .B(n5554), .Z(n5745) );
  IV U3905 ( .A(U7_DATA1_20), .Z(n5554) );
  AN2 U3906 ( .A(U7_DATA1_20), .B(n5746), .Z(n5744) );
  IV U3907 ( .A(U7_DATA1_1), .Z(n5746) );
  OR2 U3908 ( .A(n5747), .B(n5748), .Z(n5743) );
  OR2 U3909 ( .A(n279), .B(n5749), .Z(n5748) );
  AN2 U3910 ( .A(ENCODER_DATA_IN[1]), .B(n4445), .Z(n5749) );
  AN2 U3911 ( .A(U10_DATA2_1), .B(n4446), .Z(n5747) );
  AN2 U3912 ( .A(n5750), .B(n5751), .Z(ENCODER_DATA_OUT[2]) );
  IV U3913 ( .A(n5752), .Z(n5751) );
  AN2 U3914 ( .A(n5753), .B(n5754), .Z(n5752) );
  OR2 U3915 ( .A(n5754), .B(n5753), .Z(n5750) );
  OR2 U3916 ( .A(n5755), .B(n5756), .Z(n5753) );
  AN2 U3917 ( .A(U7_DATA1_0), .B(n5575), .Z(n5756) );
  IV U3918 ( .A(U7_DATA1_19), .Z(n5575) );
  AN2 U3919 ( .A(U7_DATA1_19), .B(n5757), .Z(n5755) );
  IV U3920 ( .A(U7_DATA1_0), .Z(n5757) );
  OR2 U3921 ( .A(n5758), .B(n5759), .Z(n5754) );
  OR2 U3922 ( .A(n281), .B(n5760), .Z(n5759) );
  AN2 U3923 ( .A(ENCODER_DATA_IN[0]), .B(n4445), .Z(n5760) );
  AN2 U3924 ( .A(n2491), .B(ENCODER_DATA_OUT[1]), .Z(n4445) );
  AN2 U3925 ( .A(U10_DATA2_0), .B(n4446), .Z(n5758) );
  AN2 U3926 ( .A(n2491), .B(ENCODER_DATA_OUT[0]), .Z(n4446) );
  IV U3927 ( .A(n1970), .Z(n2491) );
  IV U3928 ( .A(ENCODER_DATA_OUT[1]), .Z(ENCODER_DATA_OUT[0]) );
endmodule

