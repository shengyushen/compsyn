
module pcs_tx_dpath ( txclk, reset_tx, txd, tx_en, tx_er, adver_reg, ack, 
        txd_sel, tx_enc_ctrl_sel, tx_enc_conf_sel, link_up_loc, 
        jitter_study_pci, tx_10bdata, tx_en_d, tx_er_d, txd_eq_crs_ext, 
        pos_disp_tx_p, assertion_shengyushen );
  input [7:0] txd;
  input [12:0] adver_reg;
  input [1:0] txd_sel;
  input [3:0] tx_enc_ctrl_sel;
  input [3:0] tx_enc_conf_sel;
  input [1:0] jitter_study_pci;
  output [9:0] tx_10bdata;
  input txclk, reset_tx, tx_en, tx_er, ack, link_up_loc;
  output tx_en_d, tx_er_d, txd_eq_crs_ext, pos_disp_tx_p,
         assertion_shengyushen;
  wire   special_char, special_enc_in, pos_disp_tx, N4, N5, N6, N7, N8, N9,
         N10, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52,
         N55, N56, N57, N60, N61, N62, N65, N66, N67, N71, N72, N73, N78, N79,
         N80, N84, N85, N86, N89, N90, N91, N95, N96, N97, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N210, N1011, N911, N811, N711, N611, N511, N411, N212, N213,
         N11811, N1180, N1177, N1158, N1154, N1120, N1116, N11011, N1097,
         N1063, N1027, N9911, N976, N955, N952, N932, N922, N908, N904, N889,
         N887, N886, N885, N884, N883, N882, N8811, N870, N869, N868, N864,
         N863, N8611, N860, N859, N855, N854, N852, N850, N848, N847, N845,
         N844, N843, N842, N8411, N840, N839, N838, N837, N836, N835, N834,
         N833, N832, N8311, N830, N829, N828, N827, N826, N825, N823, N822,
         N820, N819, N817, N815, N814, N8121, N8101, N808, N806, N804, N802,
         N800, N798, N796, N794, N792, N7911, N790, N788, N787, N786, N784,
         N782, N780, N779, N777, N775, N774, N772, N7711, N769, N768, N767,
         N765, N764, N763, N7611, N760, N758, N757, N755, N754, N753, N7511,
         N750, N748, N747, N746, N745, N744, N743, N7411, N740, N739, N737,
         N736, N735, N733, N7311, N729, N727, N725, N723, N7211, N719, N717,
         N715, N7131, N7111, N709, N707, N706, N705, N703, N7011, N700, N698,
         N696, N694, N692, N690, N688, N686, N685, N683, N6811, N679, N677,
         N676, N674, N672, N670, N668, N666, N665, N663, N6611, N659, N657,
         N655, N653, N6511, N649, N647, N645, N643, N6411, N639, N637, N635,
         N633, N632, N630, N628, N626, N624, N622, N620, N618, N616, N614,
         N6121, N6101, N608, N606, N604, N602, N600, N599, N597, N595, N593,
         N5911, N589, N587, N585, N583, N5811, N579, N577, N575, N573, N5711,
         N569, N567, N566, N564, N562, N560, N558, N556, N554, N552, N550,
         N548, N546, N544, N542, N540, N538, N536, N534, N533, N532, N530,
         N528, N526, N524, N522, N520, N518, N516, N514, N5121, N5101, N508,
         N506, N504, N502, N500, N499, N498, N496, N494, N492, N490, N488,
         N486, N484, N482, N480, N478, N476, N474, N472, N470, N468, N466,
         N465, N464, N463, N4611, N459, N457, N455, N453, N4511, N449, N447,
         N445, N443, N4411, N439, N437, N435, N433, N4311, N430, N428, N426,
         N424, N422, N420, N418, N416, N414, N4121, N4101, N408, N406, N404,
         N402, N400, N398, N397, N395, N393, N3911, N389, N387, N385, N383,
         N3811, N379, N377, N375, N373, N3711, N369, N367, N365, N364, N362,
         N360, N358, N356, N354, N352, N350, N348, N346, N344, N342, N340,
         N338, N336, N334, N332, N3311, N329, N327, N326, N324, N323, N3211,
         N319, N318, N316, N3141, N3121, N3101, N308, N306, N304, N302, N300,
         N298, N296, N295, N294, N293, N2911, N290, N289, N287, N285, N283,
         N282, N280, N278, N277, N275, N274, N272, N2711, N270, N268, N267,
         N266, N264, N263, N2611, N260, N258, N257, N256, N255, N253, N252,
         N250, N249, N248, N246, N245, N244, N243, N242, N2411, N240, N239,
         N238, N237, N236, N235, N234, N233, N7061, N7051, N6971, N6721, N6701,
         N6641, N6371, N6361, N6351, N6341, N6331, N6321, N6312, N6301, N6291,
         N6281, N6271, N6261, N6251, N6241, N6231, N6221, N6212, N6201, N6191,
         N6181, N6171, N6161, N6141, N6132, N6122, N6102, N6091, N6081, N6061,
         N6041, N6031, N6012, N5991, N5971, N5951, N5941, N5931, N5912, N5891,
         N5871, N5861, N5841, N5821, N5812, N5791, N5781, N5761, N5751, N5741,
         N5731, N5721, N5701, N5691, N5681, N5671, N5651, N5631, N5612, N5601,
         N5581, N5561, N5551, N5531, N5521, N5501, N5491, N5481, N5471, N5461,
         N5451, N5441, N5421, N5401, N5391, N5371, N5361, N5341, N5321, N5312,
         N5291, N5271, N5251, N5241, N5221, N5201, N5181, N5161, N5141, N5122,
         N5102, N5081, N5061, N5051, N5041, N5021, N5001, N4981, N4961, N4941,
         N4921, N4901, N4891, N4871, N4851, N4831, N4812, N4791, N4771, N4751,
         N4741, N4721, N4701, N4681, N4661, N4651, N4631, N4612, N4591, N4571,
         N4551, N4541, N4531, N4512, N4491, N4471, N4451, N4431, N4412, N4391,
         N4371, N4351, N4331, N4312, N4291, N4271, N4251, N4231, N4212, N4201,
         N4181, N4161, N4141, N4122, N4102, N4081, N4061, N4041, N4021, N4001,
         N3981, N3961, N3941, N3921, N3901, N3881, N3871, N3851, N3831, N3812,
         N3791, N3771, N3751, N3731, N3712, N3691, N3671, N3651, N3631, N3612,
         N3591, N3571, N3561, N3541, N3521, N3501, N3481, N3461, N3441, N3421,
         N3401, N3381, N3361, N3341, N3321, N3301, N3281, N3271, N3261, N3241,
         N3221, N3201, N3181, N3161, N3142, N3122, N3102, N3081, N3061, N3041,
         N3021, N3001, N2981, N2961, N2941, N2921, N2901, N2881, N2871, N2851,
         N2831, N2812, N2791, N2771, N2751, N2731, N2712, N2691, N2671, N2651,
         N2631, N2612, N2591, N2571, N2551, N2541, N2521, N2501, N2481, N2461,
         N2441, N2421, N2401, N2381, N2361, N2341, N2321, N2301, N2281, N2261,
         N2241, N2221, N2212, N2191, N2171, N2152, N2132, N2112, N2091, N2071,
         N2051, N2031, N2012, N1991, N1971, N1951, N1931, N1912, N1891, N1881,
         N1871, N1851, N1831, N1812, N1791, N1771, N1751, N1731, N1712, N1691,
         N1671, N1651, N1631, N1612, N1591, N1571, N1551, N1541, N1531, N1512,
         N1501, N1481, N1461, N1441, N1421, N1401, N1381, N1361, N1351, N1331,
         N1312, N1291, N1271, N1251, N1231, N1212, N1192, N1187, N11710,
         N11510, N11310, N11110, N10910, N10710, N10510, N10310, N10110, N9910,
         N9710, N9510, N9310, N9210, N9010, N8810, N8710, N8510, N8410, N8310,
         N8210, N8010, N7810, N7610, N7510, N7310, N7210, N7010, N6910, N6810,
         N6610, N6510, N6310, N6210, N6010, N5910, N5810, N5610, N5410, N5310,
         N5110, N5010, N4910, N4710, N4610, N4510, N4410, N4210, N4010, N3910,
         N3810, N3710, N3610, N3510, N3310, N3110, N3010, N2910, N2810, N2710,
         N2610, N2510, N2410, N1410, N1186, rst_reg, N2103, N1190, N10102,
         N8102, N6103, N5103, N2105, sync1, sync11, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35, n37, n38,
         n40, n41, n43, n44, n48, n50, n51, n52, n53, n54, n56, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n87, n88, n89, n90, n95,
         n96, n97, n99, n100, n101, n102, n103, n105, n107, n108, n111, n112,
         n113, n114, n119, n120, n123, n124, n125, n126, n131, n132, n133,
         n135, n136, n137, n138, n139, n141, n143, n144, n145, n147, n148,
         n150, n152, n153, n154, n155, n157, n158, n161, n162, n165, n166,
         n168, n169, n172, n173, n174, n175, n176, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n195, n196, n197, n198, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n220, n221,
         n222, n223, n224, n226, n228, n229, n230, n231, n233, n234, n235,
         n236, n237, n239, n241, n242, n245, n246, n247, n248, n253, n254,
         n257, n258, n259, n260, n265, n266, n267, n269, n270, n271, n272,
         n273, n275, n277, n278, n279, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025;
  wire   [3:0] tx_enc_sel;
  wire   [7:0] txd_d;
  wire   [6:0] tx_8bdata_conf;
  wire   [7:0] tx_8b_enc_in;
  wire   [3:0] encoder_sel;
  wire   [9:0] tx_10b_enc_out;
  wire   [9:0] tx_10bdata_todiag;
  wire   [7:3] tx_10bdata_predel;
  wire   [1:0] jitter_study_tx;
  wire   [3:0] tx_enc_ctrl_sel_reg;

  IV I_09 ( .A(link_up_loc), .Z(N2105) );
  AN2 C63 ( .A(n306), .B(n308), .Z(N5103) );
  OR2 C84 ( .A(jitter_study_tx[1]), .B(n308), .Z(N6103) );
  OR2 C1113 ( .A(n306), .B(jitter_study_tx[0]), .Z(N8102) );
  AN2 C131 ( .A(jitter_study_tx[1]), .B(jitter_study_tx[0]), .Z(N10102) );
  OR2 C332 ( .A(n305), .B(N10102), .Z(N1190) );
  IV I_07 ( .A(reset_tx), .Z(N2103) );
  AN2 C272 ( .A(n289), .B(n288), .Z(N2410) );
  AN2 C282 ( .A(n287), .B(n286), .Z(N2510) );
  AN2 C292 ( .A(n285), .B(n284), .Z(N2610) );
  AN2 C303 ( .A(n283), .B(n152), .Z(N2710) );
  AN2 C312 ( .A(N2410), .B(N2510), .Z(N2810) );
  AN2 C321 ( .A(N2610), .B(N2710), .Z(N2910) );
  AN2 C331 ( .A(N2810), .B(N2910), .Z(N3010) );
  OR2 C41 ( .A(N3810), .B(N8410), .Z(N3110) );
  OR2 C502 ( .A(N3810), .B(N8710), .Z(N3310) );
  OR2 C54 ( .A(tx_8b_enc_in[7]), .B(tx_8b_enc_in[6]), .Z(N3510) );
  OR2 C551 ( .A(tx_8b_enc_in[5]), .B(tx_8b_enc_in[4]), .Z(N3610) );
  OR2 C571 ( .A(n283), .B(n152), .Z(N3710) );
  OR2 C582 ( .A(N3510), .B(N3610), .Z(N3810) );
  OR2 C591 ( .A(N5731), .B(N3710), .Z(N3910) );
  OR2 C601 ( .A(N3810), .B(N3910), .Z(N4010) );
  OR2 C692 ( .A(N3810), .B(N9210), .Z(N4210) );
  OR2 C751 ( .A(tx_8b_enc_in[3]), .B(n284), .Z(N4410) );
  OR2 C761 ( .A(tx_8b_enc_in[1]), .B(n152), .Z(N4510) );
  OR2 C781 ( .A(N4410), .B(N4510), .Z(N4610) );
  OR2 C791 ( .A(N3810), .B(N4610), .Z(N4710) );
  OR2 C86 ( .A(n283), .B(tx_8b_enc_in[0]), .Z(N4910) );
  OR2 C882 ( .A(N4410), .B(N4910), .Z(N5010) );
  OR2 C892 ( .A(N3810), .B(N5010), .Z(N5110) );
  OR2 C992 ( .A(N4410), .B(N3710), .Z(N5310) );
  OR2 C1001 ( .A(N3810), .B(N5310), .Z(N5410) );
  OR2 C1092 ( .A(N3810), .B(N1351), .Z(N5610) );
  OR2 C1151 ( .A(n285), .B(tx_8b_enc_in[2]), .Z(N5810) );
  OR2 C1182 ( .A(N5810), .B(N4510), .Z(N5910) );
  OR2 C1192 ( .A(N3810), .B(N5910), .Z(N6010) );
  OR2 C1281 ( .A(N5810), .B(N4910), .Z(N6210) );
  OR2 C129 ( .A(N3810), .B(N6210), .Z(N6310) );
  OR2 C1391 ( .A(N5810), .B(N3710), .Z(N6510) );
  OR2 C1401 ( .A(N3810), .B(N6510), .Z(N6610) );
  OR2 C146 ( .A(n285), .B(n284), .Z(N6810) );
  OR2 C149 ( .A(N6810), .B(N5471), .Z(N6910) );
  OR2 C150 ( .A(N3810), .B(N6910), .Z(N7010) );
  OR2 C160 ( .A(N6810), .B(N4510), .Z(N7210) );
  OR2 C161 ( .A(N3810), .B(N7210), .Z(N7310) );
  OR2 C1711 ( .A(N6810), .B(N4910), .Z(N7510) );
  OR2 C172 ( .A(N3810), .B(N7510), .Z(N7610) );
  OR2 C184 ( .A(N3810), .B(N1501), .Z(N7810) );
  OR2 C1931 ( .A(N8310), .B(N5751), .Z(N8010) );
  OR2 C198 ( .A(tx_8b_enc_in[5]), .B(n286), .Z(N8210) );
  OR2 C2011 ( .A(N3510), .B(N8210), .Z(N8310) );
  OR2 C202 ( .A(N5731), .B(N4510), .Z(N8410) );
  OR2 C2031 ( .A(N8310), .B(N8410), .Z(N8510) );
  OR2 C212 ( .A(N5731), .B(N4910), .Z(N8710) );
  OR2 C213 ( .A(N8310), .B(N8710), .Z(N8810) );
  OR2 C2241 ( .A(N8310), .B(N3910), .Z(N9010) );
  OR2 C233 ( .A(N4410), .B(N5471), .Z(N9210) );
  OR2 C234 ( .A(N8310), .B(N9210), .Z(N9310) );
  OR2 C245 ( .A(N8310), .B(N4610), .Z(N9510) );
  OR2 C256 ( .A(N8310), .B(N5010), .Z(N9710) );
  OR2 C2681 ( .A(N8310), .B(N5310), .Z(N9910) );
  OR2 C278 ( .A(N8310), .B(N1351), .Z(N10110) );
  OR2 C289 ( .A(N8310), .B(N5910), .Z(N10310) );
  OR2 C300 ( .A(N8310), .B(N6210), .Z(N10510) );
  OR2 C3121 ( .A(N8310), .B(N6510), .Z(N10710) );
  OR2 C323 ( .A(N8310), .B(N6910), .Z(N10910) );
  OR2 C335 ( .A(N8310), .B(N7210), .Z(N11110) );
  OR2 C347 ( .A(N8310), .B(N7510), .Z(N11310) );
  OR2 C360 ( .A(N8310), .B(N1501), .Z(N11510) );
  OR2 C364 ( .A(n287), .B(tx_8b_enc_in[4]), .Z(N11710) );
  OR2 C367 ( .A(N3510), .B(N11710), .Z(N1187) );
  OR2 C3691 ( .A(N1187), .B(N5751), .Z(N1192) );
  OR2 C3791 ( .A(N1187), .B(N8410), .Z(N1212) );
  OR2 C389 ( .A(N1187), .B(N8710), .Z(N1231) );
  OR2 C4001 ( .A(N1187), .B(N3910), .Z(N1251) );
  OR2 C410 ( .A(N1187), .B(N9210), .Z(N1271) );
  OR2 C421 ( .A(N1187), .B(N4610), .Z(N1291) );
  OR2 C432 ( .A(N1187), .B(N5010), .Z(N1312) );
  OR2 C4441 ( .A(N1187), .B(N5310), .Z(N1331) );
  OR2 C453 ( .A(N5810), .B(N5471), .Z(N1351) );
  OR2 C454 ( .A(N1187), .B(N1351), .Z(N1361) );
  OR2 C465 ( .A(N1187), .B(N5910), .Z(N1381) );
  OR2 C476 ( .A(N1187), .B(N6210), .Z(N1401) );
  OR2 C488 ( .A(N1187), .B(N6510), .Z(N1421) );
  OR2 C499 ( .A(N1187), .B(N6910), .Z(N1441) );
  OR2 C511 ( .A(N1187), .B(N7210), .Z(N1461) );
  OR2 C523 ( .A(N1187), .B(N7510), .Z(N1481) );
  OR2 C535 ( .A(N6810), .B(N3710), .Z(N1501) );
  OR2 C5361 ( .A(N1187), .B(N1501), .Z(N1512) );
  OR2 C541 ( .A(n287), .B(n286), .Z(N1531) );
  OR2 C544 ( .A(N3510), .B(N1531), .Z(N1541) );
  OR2 C546 ( .A(N1541), .B(N5751), .Z(N1551) );
  OR2 C557 ( .A(N1541), .B(N8410), .Z(N1571) );
  OR2 C568 ( .A(N1541), .B(N8710), .Z(N1591) );
  OR2 C580 ( .A(N1541), .B(N3910), .Z(N1612) );
  OR2 C5918 ( .A(N1541), .B(N9210), .Z(N1631) );
  OR2 C603 ( .A(N1541), .B(N4610), .Z(N1651) );
  OR2 C615 ( .A(N1541), .B(N5010), .Z(N1671) );
  OR2 C628 ( .A(N1541), .B(N5310), .Z(N1691) );
  OR2 C639 ( .A(N1541), .B(N1351), .Z(N1712) );
  OR2 C651 ( .A(N1541), .B(N5910), .Z(N1731) );
  OR2 C663 ( .A(N1541), .B(N6210), .Z(N1751) );
  OR2 C676 ( .A(N1541), .B(N6510), .Z(N1771) );
  OR2 C688 ( .A(N1541), .B(N6910), .Z(N1791) );
  OR2 C701 ( .A(N1541), .B(N7210), .Z(N1812) );
  OR2 C714 ( .A(N1541), .B(N7510), .Z(N1831) );
  OR2 C728 ( .A(N1541), .B(N1501), .Z(N1851) );
  OR2 C731 ( .A(tx_8b_enc_in[7]), .B(n288), .Z(N1871) );
  OR2 C735 ( .A(N1871), .B(N3610), .Z(N1881) );
  OR2 C7371 ( .A(N1881), .B(N5751), .Z(N1891) );
  OR2 C7471 ( .A(N1881), .B(N8410), .Z(N1912) );
  OR2 C757 ( .A(N1881), .B(N8710), .Z(N1931) );
  OR2 C7681 ( .A(N1881), .B(N3910), .Z(N1951) );
  OR2 C778 ( .A(N1881), .B(N9210), .Z(N1971) );
  OR2 C789 ( .A(N1881), .B(N4610), .Z(N1991) );
  OR2 C800 ( .A(N1881), .B(N5010), .Z(N2012) );
  OR2 C8121 ( .A(N1881), .B(N5310), .Z(N2031) );
  OR2 C822 ( .A(N1881), .B(N1351), .Z(N2051) );
  OR2 C833 ( .A(N1881), .B(N5910), .Z(N2071) );
  OR2 C844 ( .A(N1881), .B(N6210), .Z(N2091) );
  OR2 C856 ( .A(N1881), .B(N6510), .Z(N2112) );
  OR2 C867 ( .A(N1881), .B(N6910), .Z(N2132) );
  OR2 C879 ( .A(N1881), .B(N7210), .Z(N2152) );
  OR2 C8911 ( .A(N1881), .B(N7510), .Z(N2171) );
  OR2 C9041 ( .A(N1881), .B(N1501), .Z(N2191) );
  OR2 C912 ( .A(N1871), .B(N8210), .Z(N2212) );
  OR2 C914 ( .A(N2212), .B(N5751), .Z(N2221) );
  OR2 C925 ( .A(N2212), .B(N8410), .Z(N2241) );
  OR2 C936 ( .A(N2212), .B(N8710), .Z(N2261) );
  OR2 C948 ( .A(N2212), .B(N3910), .Z(N2281) );
  OR2 C959 ( .A(N2212), .B(N9210), .Z(N2301) );
  OR2 C971 ( .A(N2212), .B(N4610), .Z(N2321) );
  OR2 C983 ( .A(N2212), .B(N5010), .Z(N2341) );
  OR2 C996 ( .A(N2212), .B(N5310), .Z(N2361) );
  OR2 C1007 ( .A(N2212), .B(N1351), .Z(N2381) );
  OR2 C1019 ( .A(N2212), .B(N5910), .Z(N2401) );
  OR2 C1031 ( .A(N2212), .B(N6210), .Z(N2421) );
  OR2 C1044 ( .A(N2212), .B(N6510), .Z(N2441) );
  OR2 C1056 ( .A(N2212), .B(N6910), .Z(N2461) );
  OR2 C1069 ( .A(N2212), .B(N7210), .Z(N2481) );
  OR2 C1082 ( .A(N2212), .B(N7510), .Z(N2501) );
  OR2 C10961 ( .A(N2212), .B(N1501), .Z(N2521) );
  OR2 C1104 ( .A(N1871), .B(N11710), .Z(N2541) );
  OR2 C1106 ( .A(N2541), .B(N5751), .Z(N2551) );
  OR2 C1117 ( .A(N2541), .B(N8410), .Z(N2571) );
  OR2 C1128 ( .A(N2541), .B(N8710), .Z(N2591) );
  OR2 C1140 ( .A(N2541), .B(N3910), .Z(N2612) );
  OR2 C11511 ( .A(N2541), .B(N9210), .Z(N2631) );
  OR2 C1163 ( .A(N2541), .B(N4610), .Z(N2651) );
  OR2 C1175 ( .A(N2541), .B(N5010), .Z(N2671) );
  OR2 C1188 ( .A(N2541), .B(N5310), .Z(N2691) );
  OR2 C1199 ( .A(N2541), .B(N1351), .Z(N2712) );
  OR2 C1211 ( .A(N2541), .B(N5910), .Z(N2731) );
  OR2 C1223 ( .A(N2541), .B(N6210), .Z(N2751) );
  OR2 C1236 ( .A(N2541), .B(N6510), .Z(N2771) );
  OR2 C1248 ( .A(N2541), .B(N6910), .Z(N2791) );
  OR2 C1261 ( .A(N2541), .B(N7210), .Z(N2812) );
  OR2 C1274 ( .A(N2541), .B(N7510), .Z(N2831) );
  OR2 C1288 ( .A(N2541), .B(N1501), .Z(N2851) );
  OR2 C1297 ( .A(N1871), .B(N1531), .Z(N2871) );
  OR2 C1299 ( .A(N2871), .B(N5751), .Z(N2881) );
  OR2 C1311 ( .A(N2871), .B(N8410), .Z(N2901) );
  OR2 C1323 ( .A(N2871), .B(N8710), .Z(N2921) );
  OR2 C1336 ( .A(N2871), .B(N3910), .Z(N2941) );
  OR2 C1348 ( .A(N2871), .B(N9210), .Z(N2961) );
  OR2 C1361 ( .A(N2871), .B(N4610), .Z(N2981) );
  OR2 C1374 ( .A(N2871), .B(N5010), .Z(N3001) );
  OR2 C1388 ( .A(N2871), .B(N5310), .Z(N3021) );
  OR2 C1400 ( .A(N2871), .B(N1351), .Z(N3041) );
  OR2 C1413 ( .A(N2871), .B(N5910), .Z(N3061) );
  OR2 C1426 ( .A(N2871), .B(N6210), .Z(N3081) );
  OR2 C1440 ( .A(N2871), .B(N6510), .Z(N3102) );
  OR2 C1453 ( .A(N2871), .B(N6910), .Z(N3122) );
  OR2 C1467 ( .A(N2871), .B(N7210), .Z(N3142) );
  OR2 C1481 ( .A(N2871), .B(N7510), .Z(N3161) );
  OR2 C1496 ( .A(N2871), .B(N1501), .Z(N3181) );
  OR2 C15051 ( .A(N3271), .B(N5751), .Z(N3201) );
  OR2 C15151 ( .A(N3271), .B(N8410), .Z(N3221) );
  OR2 C1525 ( .A(N3271), .B(N8710), .Z(N3241) );
  OR2 C1530 ( .A(n289), .B(tx_8b_enc_in[6]), .Z(N3261) );
  OR2 C1534 ( .A(N3261), .B(N3610), .Z(N3271) );
  OR2 C15361 ( .A(N3271), .B(N3910), .Z(N3281) );
  OR2 C1546 ( .A(N3271), .B(N9210), .Z(N3301) );
  OR2 C1557 ( .A(N3271), .B(N4610), .Z(N3321) );
  OR2 C1568 ( .A(N3271), .B(N5010), .Z(N3341) );
  OR2 C15801 ( .A(N3271), .B(N5310), .Z(N3361) );
  OR2 C1590 ( .A(N3271), .B(N1351), .Z(N3381) );
  OR2 C1601 ( .A(N3271), .B(N5910), .Z(N3401) );
  OR2 C1612 ( .A(N3271), .B(N6210), .Z(N3421) );
  OR2 C1624 ( .A(N3271), .B(N6510), .Z(N3441) );
  OR2 C1635 ( .A(N3271), .B(N6910), .Z(N3461) );
  OR2 C1647 ( .A(N3271), .B(N7210), .Z(N3481) );
  OR2 C1659 ( .A(N3271), .B(N7510), .Z(N3501) );
  OR2 C16721 ( .A(N3271), .B(N1501), .Z(N3521) );
  OR2 C1682 ( .A(N3561), .B(N5751), .Z(N3541) );
  OR2 C1691 ( .A(N3261), .B(N8210), .Z(N3561) );
  OR2 C1693 ( .A(N3561), .B(N8410), .Z(N3571) );
  OR2 C1704 ( .A(N3561), .B(N8710), .Z(N3591) );
  OR2 C1716 ( .A(N3561), .B(N3910), .Z(N3612) );
  OR2 C1727 ( .A(N3561), .B(N9210), .Z(N3631) );
  OR2 C1739 ( .A(N3561), .B(N4610), .Z(N3651) );
  OR2 C1751 ( .A(N3561), .B(N5010), .Z(N3671) );
  OR2 C1764 ( .A(N3561), .B(N5310), .Z(N3691) );
  OR2 C1775 ( .A(N3561), .B(N1351), .Z(N3712) );
  OR2 C1787 ( .A(N3561), .B(N5910), .Z(N3731) );
  OR2 C1799 ( .A(N3561), .B(N6210), .Z(N3751) );
  OR2 C1812 ( .A(N3561), .B(N6510), .Z(N3771) );
  OR2 C1824 ( .A(N3561), .B(N6910), .Z(N3791) );
  OR2 C1837 ( .A(N3561), .B(N7210), .Z(N3812) );
  OR2 C1850 ( .A(N3561), .B(N7510), .Z(N3831) );
  OR2 C18641 ( .A(N3561), .B(N1501), .Z(N3851) );
  OR2 C1872 ( .A(N3261), .B(N11710), .Z(N3871) );
  OR2 C1874 ( .A(N3871), .B(N5751), .Z(N3881) );
  OR2 C1885 ( .A(N3871), .B(N8410), .Z(N3901) );
  OR2 C1896 ( .A(N3871), .B(N8710), .Z(N3921) );
  OR2 C1908 ( .A(N3871), .B(N3910), .Z(N3941) );
  OR2 C1919 ( .A(N3871), .B(N9210), .Z(N3961) );
  OR2 C19311 ( .A(N3871), .B(N4610), .Z(N3981) );
  OR2 C1943 ( .A(N3871), .B(N5010), .Z(N4001) );
  OR2 C1956 ( .A(N3871), .B(N5310), .Z(N4021) );
  OR2 C1967 ( .A(N3871), .B(N1351), .Z(N4041) );
  OR2 C1979 ( .A(N3871), .B(N5910), .Z(N4061) );
  OR2 C1991 ( .A(N3871), .B(N6210), .Z(N4081) );
  OR2 C2004 ( .A(N3871), .B(N6510), .Z(N4102) );
  OR2 C2016 ( .A(N3871), .B(N6910), .Z(N4122) );
  OR2 C2029 ( .A(N3871), .B(N7210), .Z(N4141) );
  OR2 C2042 ( .A(N3871), .B(N7510), .Z(N4161) );
  OR2 C2056 ( .A(N3871), .B(N1501), .Z(N4181) );
  OR2 C2065 ( .A(N3261), .B(N1531), .Z(N4201) );
  OR2 C2067 ( .A(N4201), .B(N5751), .Z(N4212) );
  OR2 C2079 ( .A(N4201), .B(N8410), .Z(N4231) );
  OR2 C2091 ( .A(N4201), .B(N8710), .Z(N4251) );
  OR2 C2104 ( .A(N4201), .B(N3910), .Z(N4271) );
  OR2 C2116 ( .A(N4201), .B(N9210), .Z(N4291) );
  OR2 C2129 ( .A(N4201), .B(N4610), .Z(N4312) );
  OR2 C2142 ( .A(N4201), .B(N5010), .Z(N4331) );
  OR2 C2156 ( .A(N4201), .B(N5310), .Z(N4351) );
  OR2 C2168 ( .A(N4201), .B(N1351), .Z(N4371) );
  OR2 C2181 ( .A(N4201), .B(N5910), .Z(N4391) );
  OR2 C2194 ( .A(N4201), .B(N6210), .Z(N4412) );
  OR2 C2208 ( .A(N4201), .B(N6510), .Z(N4431) );
  OR2 C2221 ( .A(N4201), .B(N6910), .Z(N4451) );
  OR2 C2235 ( .A(N4201), .B(N7210), .Z(N4471) );
  OR2 C2249 ( .A(N4201), .B(N7510), .Z(N4491) );
  OR2 C22641 ( .A(N4201), .B(N1501), .Z(N4512) );
  OR2 C2268 ( .A(n289), .B(n288), .Z(N4531) );
  OR2 C2272 ( .A(N4531), .B(N3610), .Z(N4541) );
  OR2 C2274 ( .A(N4541), .B(N5751), .Z(N4551) );
  OR2 C2285 ( .A(N4541), .B(N8410), .Z(N4571) );
  OR2 C2296 ( .A(N4541), .B(N8710), .Z(N4591) );
  OR2 C2308 ( .A(N4541), .B(N3910), .Z(N4612) );
  OR2 C2319 ( .A(N4541), .B(N9210), .Z(N4631) );
  OR2 C2330 ( .A(N4410), .B(N6081), .Z(N4651) );
  OR2 C2331 ( .A(N4541), .B(N4651), .Z(N4661) );
  OR2 C2343 ( .A(N4541), .B(N5391), .Z(N4681) );
  OR2 C2356 ( .A(N4541), .B(N5941), .Z(N4701) );
  OR2 C2367 ( .A(N4541), .B(N1351), .Z(N4721) );
  OR2 C2378 ( .A(N5810), .B(N6081), .Z(N4741) );
  OR2 C2379 ( .A(N4541), .B(N4741), .Z(N4751) );
  OR2 C2391 ( .A(N4541), .B(N5551), .Z(N4771) );
  OR2 C2404 ( .A(N4541), .B(N6031), .Z(N4791) );
  OR2 C2416 ( .A(N4541), .B(N5601), .Z(N4812) );
  OR2 C2429 ( .A(N4541), .B(N6091), .Z(N4831) );
  OR2 C2442 ( .A(N4541), .B(N6132), .Z(N4851) );
  OR2 C2456 ( .A(N4541), .B(N5691), .Z(N4871) );
  OR2 C2465 ( .A(N4531), .B(N8210), .Z(N4891) );
  OR2 C2467 ( .A(N4891), .B(N5751), .Z(N4901) );
  OR2 C24791 ( .A(N4891), .B(N5781), .Z(N4921) );
  OR2 C2491 ( .A(N5051), .B(N5812), .Z(N4941) );
  OR2 C2504 ( .A(N5051), .B(N5312), .Z(N4961) );
  OR2 C2516 ( .A(N5051), .B(N5861), .Z(N4981) );
  OR2 C2529 ( .A(N5051), .B(N5361), .Z(N5001) );
  OR2 C2542 ( .A(N5051), .B(N5391), .Z(N5021) );
  OR2 C2551 ( .A(tx_8b_enc_in[5]), .B(n286), .Z(N5041) );
  OR2 C2554 ( .A(N4531), .B(N5041), .Z(N5051) );
  OR2 C2556 ( .A(N5051), .B(N5941), .Z(N5061) );
  OR2 C2568 ( .A(N5051), .B(N5491), .Z(N5081) );
  OR2 C2581 ( .A(N5051), .B(N5521), .Z(N5102) );
  OR2 C2594 ( .A(N5051), .B(N5551), .Z(N5122) );
  OR2 C2608 ( .A(N5051), .B(N6031), .Z(N5141) );
  OR2 C2621 ( .A(N5051), .B(N5601), .Z(N5161) );
  OR2 C2635 ( .A(N5051), .B(N6091), .Z(N5181) );
  OR2 C2649 ( .A(N5051), .B(N6132), .Z(N5201) );
  OR2 C2664 ( .A(N5051), .B(N5691), .Z(N5221) );
  OR2 C2673 ( .A(N4531), .B(N11710), .Z(N5241) );
  OR2 C2675 ( .A(N5241), .B(N5751), .Z(N5251) );
  OR2 C26871 ( .A(N5241), .B(N5781), .Z(N5271) );
  OR2 C2699 ( .A(N5481), .B(N5812), .Z(N5291) );
  OR2 C2711 ( .A(N5731), .B(N5681), .Z(N5312) );
  OR2 C2712 ( .A(N5481), .B(N5312), .Z(N5321) );
  OR2 C2724 ( .A(N5481), .B(N5861), .Z(N5341) );
  OR2 C2736 ( .A(N5931), .B(N6081), .Z(N5361) );
  OR2 C2737 ( .A(N5481), .B(N5361), .Z(N5371) );
  OR2 C2749 ( .A(N5931), .B(N6122), .Z(N5391) );
  OR2 C2750 ( .A(N5481), .B(N5391), .Z(N5401) );
  OR2 C2764 ( .A(N5481), .B(N5941), .Z(N5421) );
  OR2 C2770 ( .A(n289), .B(n288), .Z(N5441) );
  OR2 C2771 ( .A(n287), .B(tx_8b_enc_in[4]), .Z(N5451) );
  OR2 C2772 ( .A(n285), .B(tx_8b_enc_in[2]), .Z(N5461) );
  OR2 C2773 ( .A(tx_8b_enc_in[1]), .B(tx_8b_enc_in[0]), .Z(N5471) );
  OR2 C2774 ( .A(N5441), .B(N5451), .Z(N5481) );
  OR2 C2775 ( .A(N5461), .B(N5471), .Z(N5491) );
  OR2 C2776 ( .A(N5481), .B(N5491), .Z(N5501) );
  OR2 C2788 ( .A(N5461), .B(N6081), .Z(N5521) );
  OR2 C2789 ( .A(N5481), .B(N5521), .Z(N5531) );
  OR2 C2801 ( .A(N5461), .B(N6122), .Z(N5551) );
  OR2 C2802 ( .A(N5481), .B(N5551), .Z(N5561) );
  OR2 C2816 ( .A(N5481), .B(N6031), .Z(N5581) );
  OR2 C2828 ( .A(N5671), .B(N5471), .Z(N5601) );
  OR2 C2829 ( .A(N5481), .B(N5601), .Z(N5612) );
  OR2 C2843 ( .A(N5481), .B(N6091), .Z(N5631) );
  OR2 C2857 ( .A(N5481), .B(N6132), .Z(N5651) );
  OR2 C2868 ( .A(n285), .B(n284), .Z(N5671) );
  OR2 C28691 ( .A(n283), .B(n152), .Z(N5681) );
  OR2 C2871 ( .A(N5671), .B(N5681), .Z(N5691) );
  OR2 C28721 ( .A(N5481), .B(N5691), .Z(N5701) );
  OR2 C2879 ( .A(n287), .B(n286), .Z(N5721) );
  OR2 C2880 ( .A(tx_8b_enc_in[3]), .B(tx_8b_enc_in[2]), .Z(N5731) );
  OR2 C2882 ( .A(N5441), .B(N5721), .Z(N5741) );
  OR2 C2883 ( .A(N5731), .B(N5471), .Z(N5751) );
  OR2 C2884 ( .A(N5741), .B(N5751), .Z(N5761) );
  OR2 C2896 ( .A(N5731), .B(N6081), .Z(N5781) );
  OR2 C2897 ( .A(N5741), .B(N5781), .Z(N5791) );
  OR2 C2909 ( .A(N5731), .B(N6122), .Z(N5812) );
  OR2 C2910 ( .A(N5741), .B(N5812), .Z(N5821) );
  OR2 C2924 ( .A(N5741), .B(N5312), .Z(N5841) );
  OR2 C2936 ( .A(N5931), .B(N5471), .Z(N5861) );
  OR2 C2937 ( .A(N5741), .B(N5861), .Z(N5871) );
  OR2 C2951 ( .A(N5741), .B(N5361), .Z(N5891) );
  OR2 C2965 ( .A(N5741), .B(N5391), .Z(N5912) );
  OR2 C2976 ( .A(tx_8b_enc_in[3]), .B(n284), .Z(N5931) );
  OR2 C2979 ( .A(N5931), .B(N5681), .Z(N5941) );
  OR2 C2980 ( .A(N5741), .B(N5941), .Z(N5951) );
  OR2 C2993 ( .A(N5741), .B(N5491), .Z(N5971) );
  OR2 C3007 ( .A(N5741), .B(N5521), .Z(N5991) );
  OR2 C3021 ( .A(N5741), .B(N5551), .Z(N6012) );
  OR2 C3035 ( .A(N5461), .B(N5681), .Z(N6031) );
  OR2 C3036 ( .A(N5741), .B(N6031), .Z(N6041) );
  OR2 C3050 ( .A(N5741), .B(N5601), .Z(N6061) );
  OR2 C3062 ( .A(tx_8b_enc_in[1]), .B(n152), .Z(N6081) );
  OR2 C3064 ( .A(N5671), .B(N6081), .Z(N6091) );
  OR2 C3065 ( .A(N5741), .B(N6091), .Z(N6102) );
  OR2 C30771 ( .A(n283), .B(tx_8b_enc_in[0]), .Z(N6122) );
  OR2 C3079 ( .A(N5671), .B(N6122), .Z(N6132) );
  OR2 C3080 ( .A(N5741), .B(N6132), .Z(N6141) );
  AN2 C3082 ( .A(tx_8b_enc_in[7]), .B(tx_8b_enc_in[6]), .Z(N6161) );
  AN2 C3083 ( .A(tx_8b_enc_in[5]), .B(tx_8b_enc_in[4]), .Z(N6171) );
  AN2 C3084 ( .A(tx_8b_enc_in[3]), .B(tx_8b_enc_in[2]), .Z(N6181) );
  AN2 C3085 ( .A(tx_8b_enc_in[1]), .B(tx_8b_enc_in[0]), .Z(N6191) );
  AN2 C3086 ( .A(N6161), .B(N6171), .Z(N6201) );
  AN2 C3087 ( .A(N6181), .B(N6191), .Z(N6212) );
  AN2 C3088 ( .A(N6201), .B(N6212), .Z(N6221) );
  OR2 C3636 ( .A(N6361), .B(N6312), .Z(N6371) );
  OR2 C3670 ( .A(n150), .B(N6641), .Z(N6701) );
  OR2 C3672 ( .A(n148), .B(N6701), .Z(N6721) );
  OR2 C3697 ( .A(n281), .B(n282), .Z(N6971) );
  AN2 C3716 ( .A(n303), .B(n302), .Z(N1186) );
  AN2 C3720 ( .A(encoder_sel[2]), .B(n301), .Z(N1410) );
  AN2 C4250 ( .A(N7051), .B(n296), .Z(N6241) );
  AN2 C4251 ( .A(N1186), .B(n301), .Z(N7051) );
  AN2 C4252 ( .A(N1186), .B(encoder_sel[0]), .Z(N6251) );
  AN2 C4253 ( .A(n302), .B(encoder_sel[1]), .Z(N6261) );
  AN2 C4254 ( .A(N1410), .B(n296), .Z(N6271) );
  AN2 C4255 ( .A(N1410), .B(encoder_sel[0]), .Z(N6281) );
  AN2 C4256 ( .A(N7061), .B(n296), .Z(N6291) );
  AN2 C4257 ( .A(encoder_sel[2]), .B(encoder_sel[1]), .Z(N7061) );
  AN2 C4258 ( .A(encoder_sel[1]), .B(encoder_sel[0]), .Z(N6301) );
  AN2 C4259 ( .A(encoder_sel[3]), .B(n296), .Z(N6312) );
  AN2 C4260 ( .A(encoder_sel[3]), .B(encoder_sel[0]), .Z(N6321) );
  AN2 C171 ( .A(n289), .B(n288), .Z(N233) );
  AN2 C182 ( .A(n287), .B(n286), .Z(N234) );
  AN2 C191 ( .A(n285), .B(n284), .Z(N235) );
  AN2 C201 ( .A(n283), .B(n152), .Z(N236) );
  AN2 C21 ( .A(N233), .B(N234), .Z(N237) );
  AN2 C22 ( .A(N235), .B(N236), .Z(N238) );
  AN2 C231 ( .A(N237), .B(N238), .Z(N239) );
  OR2 C251 ( .A(tx_8b_enc_in[7]), .B(tx_8b_enc_in[6]), .Z(N240) );
  OR2 C26 ( .A(tx_8b_enc_in[5]), .B(tx_8b_enc_in[4]), .Z(N2411) );
  OR2 C271 ( .A(tx_8b_enc_in[3]), .B(tx_8b_enc_in[2]), .Z(N242) );
  OR2 C281 ( .A(tx_8b_enc_in[1]), .B(n152), .Z(N243) );
  OR2 C291 ( .A(N240), .B(N2411), .Z(N244) );
  OR2 C30 ( .A(N242), .B(N243), .Z(N245) );
  OR2 C311 ( .A(N244), .B(N245), .Z(N246) );
  OR2 C37 ( .A(n283), .B(tx_8b_enc_in[0]), .Z(N248) );
  OR2 C391 ( .A(N242), .B(N248), .Z(N249) );
  OR2 C401 ( .A(N244), .B(N249), .Z(N250) );
  OR2 C491 ( .A(N242), .B(N266), .Z(N252) );
  OR2 C501 ( .A(N244), .B(N252), .Z(N253) );
  OR2 C55 ( .A(tx_8b_enc_in[3]), .B(n284), .Z(N255) );
  OR2 C561 ( .A(tx_8b_enc_in[1]), .B(tx_8b_enc_in[0]), .Z(N256) );
  OR2 C581 ( .A(N255), .B(N256), .Z(N257) );
  OR2 C59 ( .A(N244), .B(N257), .Z(N258) );
  OR2 C68 ( .A(N255), .B(N243), .Z(N260) );
  OR2 C69 ( .A(N244), .B(N260), .Z(N2611) );
  OR2 C78 ( .A(N255), .B(N248), .Z(N263) );
  OR2 C79 ( .A(N244), .B(N263), .Z(N264) );
  OR2 C87 ( .A(n283), .B(n152), .Z(N266) );
  OR2 C891 ( .A(N255), .B(N266), .Z(N267) );
  OR2 C901 ( .A(N244), .B(N267), .Z(N268) );
  OR2 C951 ( .A(n285), .B(tx_8b_enc_in[2]), .Z(N270) );
  OR2 C98 ( .A(N270), .B(N256), .Z(N2711) );
  OR2 C991 ( .A(N244), .B(N2711), .Z(N272) );
  OR2 C108 ( .A(N270), .B(N243), .Z(N274) );
  OR2 C109 ( .A(N244), .B(N274), .Z(N275) );
  OR2 C1181 ( .A(N270), .B(N248), .Z(N277) );
  OR2 C1191 ( .A(N244), .B(N277), .Z(N278) );
  OR2 C130 ( .A(N244), .B(N318), .Z(N280) );
  OR2 C139 ( .A(N289), .B(N256), .Z(N282) );
  OR2 C140 ( .A(N244), .B(N282), .Z(N283) );
  OR2 C151 ( .A(N244), .B(N323), .Z(N285) );
  OR2 C162 ( .A(N244), .B(N326), .Z(N287) );
  OR2 C170 ( .A(n285), .B(n284), .Z(N289) );
  OR2 C173 ( .A(N289), .B(N266), .Z(N290) );
  OR2 C174 ( .A(N244), .B(N290), .Z(N2911) );
  OR2 C178 ( .A(tx_8b_enc_in[5]), .B(n286), .Z(N293) );
  OR2 C1811 ( .A(N240), .B(N293), .Z(N294) );
  OR2 C1821 ( .A(N242), .B(N256), .Z(N295) );
  OR2 C183 ( .A(N294), .B(N295), .Z(N296) );
  OR2 C193 ( .A(N294), .B(N245), .Z(N298) );
  OR2 C203 ( .A(N294), .B(N249), .Z(N300) );
  OR2 C214 ( .A(N294), .B(N252), .Z(N302) );
  OR2 C224 ( .A(N294), .B(N257), .Z(N304) );
  OR2 C235 ( .A(N294), .B(N260), .Z(N306) );
  OR2 C246 ( .A(N294), .B(N263), .Z(N308) );
  OR2 C258 ( .A(N294), .B(N267), .Z(N3101) );
  OR2 C268 ( .A(N294), .B(N2711), .Z(N3121) );
  OR2 C279 ( .A(N294), .B(N274), .Z(N3141) );
  OR2 C290 ( .A(N294), .B(N277), .Z(N316) );
  OR2 C301 ( .A(N270), .B(N266), .Z(N318) );
  OR2 C302 ( .A(N294), .B(N318), .Z(N319) );
  OR2 C313 ( .A(N294), .B(N282), .Z(N3211) );
  OR2 C324 ( .A(N289), .B(N243), .Z(N323) );
  OR2 C325 ( .A(N294), .B(N323), .Z(N324) );
  OR2 C336 ( .A(N289), .B(N248), .Z(N326) );
  OR2 C337 ( .A(N294), .B(N326), .Z(N327) );
  OR2 C350 ( .A(N294), .B(N290), .Z(N329) );
  OR2 C357 ( .A(N240), .B(N464), .Z(N3311) );
  OR2 C359 ( .A(N3311), .B(N295), .Z(N332) );
  OR2 C369 ( .A(N3311), .B(N245), .Z(N334) );
  OR2 C379 ( .A(N3311), .B(N249), .Z(N336) );
  OR2 C390 ( .A(N3311), .B(N252), .Z(N338) );
  OR2 C400 ( .A(N3311), .B(N257), .Z(N340) );
  OR2 C411 ( .A(N3311), .B(N260), .Z(N342) );
  OR2 C422 ( .A(N3311), .B(N263), .Z(N344) );
  OR2 C434 ( .A(N3311), .B(N267), .Z(N346) );
  OR2 C444 ( .A(N3311), .B(N2711), .Z(N348) );
  OR2 C455 ( .A(N3311), .B(N274), .Z(N350) );
  OR2 C466 ( .A(N3311), .B(N277), .Z(N352) );
  OR2 C478 ( .A(N3311), .B(N318), .Z(N354) );
  OR2 C489 ( .A(N3311), .B(N282), .Z(N356) );
  OR2 C5011 ( .A(N3311), .B(N323), .Z(N358) );
  OR2 C513 ( .A(N3311), .B(N326), .Z(N360) );
  OR2 C526 ( .A(N3311), .B(N290), .Z(N362) );
  OR2 C534 ( .A(N240), .B(N498), .Z(N364) );
  OR2 C536 ( .A(N364), .B(N295), .Z(N365) );
  OR2 C547 ( .A(N364), .B(N245), .Z(N367) );
  OR2 C558 ( .A(N364), .B(N249), .Z(N369) );
  OR2 C570 ( .A(N364), .B(N252), .Z(N3711) );
  OR2 C5811 ( .A(N364), .B(N257), .Z(N373) );
  OR2 C593 ( .A(N364), .B(N260), .Z(N375) );
  OR2 C605 ( .A(N364), .B(N263), .Z(N377) );
  OR2 C618 ( .A(N364), .B(N267), .Z(N379) );
  OR2 C629 ( .A(N364), .B(N2711), .Z(N3811) );
  OR2 C641 ( .A(N364), .B(N274), .Z(N383) );
  OR2 C653 ( .A(N364), .B(N277), .Z(N385) );
  OR2 C666 ( .A(N364), .B(N318), .Z(N387) );
  OR2 C678 ( .A(N364), .B(N282), .Z(N389) );
  OR2 C691 ( .A(N364), .B(N323), .Z(N3911) );
  OR2 C704 ( .A(N364), .B(N326), .Z(N393) );
  OR2 C718 ( .A(N364), .B(N290), .Z(N395) );
  OR2 C725 ( .A(N463), .B(N2411), .Z(N397) );
  OR2 C727 ( .A(N397), .B(N295), .Z(N398) );
  OR2 C737 ( .A(N397), .B(N245), .Z(N400) );
  OR2 C747 ( .A(N397), .B(N249), .Z(N402) );
  OR2 C758 ( .A(N397), .B(N252), .Z(N404) );
  OR2 C768 ( .A(N397), .B(N257), .Z(N406) );
  OR2 C779 ( .A(N397), .B(N260), .Z(N408) );
  OR2 C790 ( .A(N397), .B(N263), .Z(N4101) );
  OR2 C802 ( .A(N397), .B(N267), .Z(N4121) );
  OR2 C812 ( .A(N397), .B(N2711), .Z(N414) );
  OR2 C823 ( .A(N397), .B(N274), .Z(N416) );
  OR2 C834 ( .A(N397), .B(N277), .Z(N418) );
  OR2 C846 ( .A(N397), .B(N318), .Z(N420) );
  OR2 C857 ( .A(N397), .B(N282), .Z(N422) );
  OR2 C869 ( .A(N397), .B(N323), .Z(N424) );
  OR2 C881 ( .A(N397), .B(N326), .Z(N426) );
  OR2 C894 ( .A(N397), .B(N290), .Z(N428) );
  OR2 C902 ( .A(N463), .B(N293), .Z(N430) );
  OR2 C904 ( .A(N430), .B(N295), .Z(N4311) );
  OR2 C915 ( .A(N430), .B(N245), .Z(N433) );
  OR2 C926 ( .A(N430), .B(N249), .Z(N435) );
  OR2 C938 ( .A(N430), .B(N252), .Z(N437) );
  OR2 C949 ( .A(N430), .B(N257), .Z(N439) );
  OR2 C961 ( .A(N430), .B(N260), .Z(N4411) );
  OR2 C973 ( .A(N430), .B(N263), .Z(N443) );
  OR2 C986 ( .A(N430), .B(N267), .Z(N445) );
  OR2 C997 ( .A(N430), .B(N2711), .Z(N447) );
  OR2 C1009 ( .A(N430), .B(N274), .Z(N449) );
  OR2 C1021 ( .A(N430), .B(N277), .Z(N4511) );
  OR2 C1034 ( .A(N430), .B(N318), .Z(N453) );
  OR2 C1046 ( .A(N430), .B(N282), .Z(N455) );
  OR2 C1059 ( .A(N430), .B(N323), .Z(N457) );
  OR2 C1072 ( .A(N430), .B(N326), .Z(N459) );
  OR2 C1086 ( .A(N430), .B(N290), .Z(N4611) );
  OR2 C1090 ( .A(tx_8b_enc_in[7]), .B(n288), .Z(N463) );
  OR2 C1091 ( .A(n287), .B(tx_8b_enc_in[4]), .Z(N464) );
  OR2 C1094 ( .A(N463), .B(N464), .Z(N465) );
  OR2 C1096 ( .A(N465), .B(N295), .Z(N466) );
  OR2 C1107 ( .A(N465), .B(N245), .Z(N468) );
  OR2 C1118 ( .A(N465), .B(N249), .Z(N470) );
  OR2 C1130 ( .A(N465), .B(N252), .Z(N472) );
  OR2 C1141 ( .A(N465), .B(N257), .Z(N474) );
  OR2 C1153 ( .A(N465), .B(N260), .Z(N476) );
  OR2 C1165 ( .A(N465), .B(N263), .Z(N478) );
  OR2 C1178 ( .A(N465), .B(N267), .Z(N480) );
  OR2 C1189 ( .A(N465), .B(N2711), .Z(N482) );
  OR2 C1201 ( .A(N465), .B(N274), .Z(N484) );
  OR2 C1213 ( .A(N465), .B(N277), .Z(N486) );
  OR2 C1226 ( .A(N465), .B(N318), .Z(N488) );
  OR2 C1238 ( .A(N465), .B(N282), .Z(N490) );
  OR2 C1251 ( .A(N465), .B(N323), .Z(N492) );
  OR2 C1264 ( .A(N465), .B(N326), .Z(N494) );
  OR2 C1278 ( .A(N465), .B(N290), .Z(N496) );
  OR2 C1284 ( .A(n287), .B(n286), .Z(N498) );
  OR2 C1287 ( .A(N463), .B(N498), .Z(N499) );
  OR2 C1289 ( .A(N499), .B(N295), .Z(N500) );
  OR2 C1301 ( .A(N499), .B(N245), .Z(N502) );
  OR2 C1313 ( .A(N499), .B(N249), .Z(N504) );
  OR2 C1326 ( .A(N499), .B(N252), .Z(N506) );
  OR2 C1338 ( .A(N499), .B(N257), .Z(N508) );
  OR2 C1351 ( .A(N499), .B(N260), .Z(N5101) );
  OR2 C1364 ( .A(N499), .B(N263), .Z(N5121) );
  OR2 C1378 ( .A(N499), .B(N267), .Z(N514) );
  OR2 C1390 ( .A(N499), .B(N2711), .Z(N516) );
  OR2 C1403 ( .A(N499), .B(N274), .Z(N518) );
  OR2 C1416 ( .A(N499), .B(N277), .Z(N520) );
  OR2 C1430 ( .A(N499), .B(N318), .Z(N522) );
  OR2 C1443 ( .A(N499), .B(N282), .Z(N524) );
  OR2 C1457 ( .A(N499), .B(N323), .Z(N526) );
  OR2 C1471 ( .A(N499), .B(N326), .Z(N528) );
  OR2 C1486 ( .A(N499), .B(N290), .Z(N530) );
  OR2 C1489 ( .A(n289), .B(tx_8b_enc_in[6]), .Z(N532) );
  OR2 C1493 ( .A(N532), .B(N2411), .Z(N533) );
  OR2 C1495 ( .A(N533), .B(N295), .Z(N534) );
  OR2 C1505 ( .A(N533), .B(N245), .Z(N536) );
  OR2 C1515 ( .A(N533), .B(N249), .Z(N538) );
  OR2 C1526 ( .A(N533), .B(N252), .Z(N540) );
  OR2 C1536 ( .A(N533), .B(N257), .Z(N542) );
  OR2 C1547 ( .A(N533), .B(N260), .Z(N544) );
  OR2 C1558 ( .A(N533), .B(N263), .Z(N546) );
  OR2 C1570 ( .A(N533), .B(N267), .Z(N548) );
  OR2 C1580 ( .A(N533), .B(N2711), .Z(N550) );
  OR2 C1591 ( .A(N533), .B(N274), .Z(N552) );
  OR2 C1602 ( .A(N533), .B(N277), .Z(N554) );
  OR2 C1614 ( .A(N533), .B(N318), .Z(N556) );
  OR2 C1625 ( .A(N533), .B(N282), .Z(N558) );
  OR2 C1637 ( .A(N533), .B(N323), .Z(N560) );
  OR2 C1649 ( .A(N533), .B(N326), .Z(N562) );
  OR2 C1662 ( .A(N533), .B(N290), .Z(N564) );
  OR2 C1670 ( .A(N532), .B(N293), .Z(N566) );
  OR2 C1672 ( .A(N566), .B(N295), .Z(N567) );
  OR2 C1683 ( .A(N566), .B(N245), .Z(N569) );
  OR2 C1694 ( .A(N566), .B(N249), .Z(N5711) );
  OR2 C1706 ( .A(N566), .B(N252), .Z(N573) );
  OR2 C1717 ( .A(N566), .B(N257), .Z(N575) );
  OR2 C1729 ( .A(N566), .B(N260), .Z(N577) );
  OR2 C1741 ( .A(N566), .B(N263), .Z(N579) );
  OR2 C1754 ( .A(N566), .B(N267), .Z(N5811) );
  OR2 C1765 ( .A(N566), .B(N2711), .Z(N583) );
  OR2 C1777 ( .A(N566), .B(N274), .Z(N585) );
  OR2 C1789 ( .A(N566), .B(N277), .Z(N587) );
  OR2 C1802 ( .A(N566), .B(N318), .Z(N589) );
  OR2 C1814 ( .A(N566), .B(N282), .Z(N5911) );
  OR2 C1827 ( .A(N566), .B(N323), .Z(N593) );
  OR2 C1840 ( .A(N566), .B(N326), .Z(N595) );
  OR2 C1854 ( .A(N566), .B(N290), .Z(N597) );
  OR2 C1862 ( .A(N532), .B(N464), .Z(N599) );
  OR2 C1864 ( .A(N599), .B(N295), .Z(N600) );
  OR2 C1875 ( .A(N599), .B(N245), .Z(N602) );
  OR2 C1886 ( .A(N599), .B(N249), .Z(N604) );
  OR2 C1898 ( .A(N599), .B(N252), .Z(N606) );
  OR2 C1909 ( .A(N599), .B(N257), .Z(N608) );
  OR2 C1921 ( .A(N599), .B(N260), .Z(N6101) );
  OR2 C1933 ( .A(N599), .B(N263), .Z(N6121) );
  OR2 C1946 ( .A(N599), .B(N267), .Z(N614) );
  OR2 C1957 ( .A(N599), .B(N2711), .Z(N616) );
  OR2 C1969 ( .A(N599), .B(N274), .Z(N618) );
  OR2 C1981 ( .A(N599), .B(N277), .Z(N620) );
  OR2 C1994 ( .A(N599), .B(N318), .Z(N622) );
  OR2 C2006 ( .A(N599), .B(N282), .Z(N624) );
  OR2 C2019 ( .A(N599), .B(N323), .Z(N626) );
  OR2 C2032 ( .A(N599), .B(N326), .Z(N628) );
  OR2 C2046 ( .A(N599), .B(N290), .Z(N630) );
  OR2 C2055 ( .A(N532), .B(N498), .Z(N632) );
  OR2 C2057 ( .A(N632), .B(N295), .Z(N633) );
  OR2 C2069 ( .A(N632), .B(N245), .Z(N635) );
  OR2 C2081 ( .A(N632), .B(N249), .Z(N637) );
  OR2 C2094 ( .A(N632), .B(N252), .Z(N639) );
  OR2 C2106 ( .A(N632), .B(N257), .Z(N6411) );
  OR2 C2119 ( .A(N632), .B(N260), .Z(N643) );
  OR2 C2132 ( .A(N632), .B(N263), .Z(N645) );
  OR2 C2146 ( .A(N632), .B(N267), .Z(N647) );
  OR2 C2158 ( .A(N632), .B(N2711), .Z(N649) );
  OR2 C2171 ( .A(N632), .B(N274), .Z(N6511) );
  OR2 C2184 ( .A(N632), .B(N277), .Z(N653) );
  OR2 C2198 ( .A(N632), .B(N318), .Z(N655) );
  OR2 C2211 ( .A(N632), .B(N282), .Z(N657) );
  OR2 C2225 ( .A(N632), .B(N323), .Z(N659) );
  OR2 C2239 ( .A(N632), .B(N326), .Z(N6611) );
  OR2 C2254 ( .A(N632), .B(N290), .Z(N663) );
  OR2 C2262 ( .A(N735), .B(N2411), .Z(N665) );
  OR2 C2264 ( .A(N665), .B(N295), .Z(N666) );
  OR2 C2275 ( .A(N665), .B(N245), .Z(N668) );
  OR2 C2286 ( .A(N665), .B(N249), .Z(N670) );
  OR2 C2298 ( .A(N665), .B(N252), .Z(N672) );
  OR2 C2309 ( .A(N665), .B(N257), .Z(N674) );
  OR2 C2320 ( .A(N255), .B(N739), .Z(N676) );
  OR2 C2321 ( .A(N665), .B(N676), .Z(N677) );
  OR2 C2333 ( .A(N665), .B(N760), .Z(N679) );
  OR2 C2346 ( .A(N665), .B(N764), .Z(N6811) );
  OR2 C2357 ( .A(N665), .B(N2711), .Z(N683) );
  OR2 C2368 ( .A(N270), .B(N739), .Z(N685) );
  OR2 C2369 ( .A(N665), .B(N685), .Z(N686) );
  OR2 C2381 ( .A(N665), .B(N774), .Z(N688) );
  OR2 C2394 ( .A(N665), .B(N814), .Z(N690) );
  OR2 C2406 ( .A(N665), .B(N779), .Z(N692) );
  OR2 C2419 ( .A(N665), .B(N819), .Z(N694) );
  OR2 C2432 ( .A(N665), .B(N822), .Z(N696) );
  OR2 C2446 ( .A(N665), .B(N787), .Z(N698) );
  OR2 C2455 ( .A(N735), .B(N293), .Z(N700) );
  OR2 C2457 ( .A(N700), .B(N295), .Z(N7011) );
  OR2 C2469 ( .A(N700), .B(N740), .Z(N703) );
  OR2 C2476 ( .A(tx_8b_enc_in[5]), .B(n286), .Z(N705) );
  OR2 C2479 ( .A(N735), .B(N705), .Z(N706) );
  OR2 C2481 ( .A(N706), .B(N747), .Z(N707) );
  OR2 C2494 ( .A(N706), .B(N750), .Z(N709) );
  OR2 C2506 ( .A(N706), .B(N754), .Z(N7111) );
  OR2 C2519 ( .A(N706), .B(N757), .Z(N7131) );
  OR2 C2532 ( .A(N706), .B(N760), .Z(N715) );
  OR2 C2546 ( .A(N706), .B(N764), .Z(N717) );
  OR2 C2558 ( .A(N706), .B(N768), .Z(N719) );
  OR2 C2571 ( .A(N706), .B(N7711), .Z(N7211) );
  OR2 C2584 ( .A(N706), .B(N774), .Z(N723) );
  OR2 C2598 ( .A(N706), .B(N814), .Z(N725) );
  OR2 C2611 ( .A(N706), .B(N779), .Z(N727) );
  OR2 C2625 ( .A(N706), .B(N819), .Z(N729) );
  OR2 C2639 ( .A(N706), .B(N822), .Z(N7311) );
  OR2 C2654 ( .A(N706), .B(N787), .Z(N733) );
  OR2 C2659 ( .A(n289), .B(n288), .Z(N735) );
  OR2 C2663 ( .A(N735), .B(N464), .Z(N736) );
  OR2 C2665 ( .A(N736), .B(N295), .Z(N737) );
  OR2 C2674 ( .A(tx_8b_enc_in[1]), .B(n152), .Z(N739) );
  OR2 C2676 ( .A(N242), .B(N739), .Z(N740) );
  OR2 C2677 ( .A(N736), .B(N740), .Z(N7411) );
  OR2 C2683 ( .A(n289), .B(n288), .Z(N743) );
  OR2 C2684 ( .A(n287), .B(tx_8b_enc_in[4]), .Z(N744) );
  OR2 C2686 ( .A(n283), .B(tx_8b_enc_in[0]), .Z(N745) );
  OR2 C2687 ( .A(N743), .B(N744), .Z(N746) );
  OR2 C2688 ( .A(N242), .B(N745), .Z(N747) );
  OR2 C2689 ( .A(N746), .B(N747), .Z(N748) );
  OR2 C2701 ( .A(N242), .B(N763), .Z(N750) );
  OR2 C2702 ( .A(N746), .B(N750), .Z(N7511) );
  OR2 C2710 ( .A(tx_8b_enc_in[3]), .B(n284), .Z(N753) );
  OR2 C2713 ( .A(N753), .B(N256), .Z(N754) );
  OR2 C2714 ( .A(N746), .B(N754), .Z(N755) );
  OR2 C2726 ( .A(N753), .B(N739), .Z(N757) );
  OR2 C2727 ( .A(N746), .B(N757), .Z(N758) );
  OR2 C2739 ( .A(N753), .B(N745), .Z(N760) );
  OR2 C2740 ( .A(N746), .B(N760), .Z(N7611) );
  OR2 C2751 ( .A(n283), .B(n152), .Z(N763) );
  OR2 C2753 ( .A(N753), .B(N763), .Z(N764) );
  OR2 C2754 ( .A(N746), .B(N764), .Z(N765) );
  OR2 C2762 ( .A(n285), .B(tx_8b_enc_in[2]), .Z(N767) );
  OR2 C2765 ( .A(N767), .B(N256), .Z(N768) );
  OR2 C2766 ( .A(N746), .B(N768), .Z(N769) );
  OR2 C2778 ( .A(N767), .B(N739), .Z(N7711) );
  OR2 C2779 ( .A(N746), .B(N7711), .Z(N772) );
  OR2 C2791 ( .A(N767), .B(N745), .Z(N774) );
  OR2 C2792 ( .A(N746), .B(N774), .Z(N775) );
  OR2 C2806 ( .A(N746), .B(N814), .Z(N777) );
  OR2 C2818 ( .A(N786), .B(N256), .Z(N779) );
  OR2 C2819 ( .A(N746), .B(N779), .Z(N780) );
  OR2 C2833 ( .A(N746), .B(N819), .Z(N782) );
  OR2 C2847 ( .A(N746), .B(N822), .Z(N784) );
  OR2 C2858 ( .A(n285), .B(n284), .Z(N786) );
  OR2 C2861 ( .A(N786), .B(N763), .Z(N787) );
  OR2 C2862 ( .A(N746), .B(N787), .Z(N788) );
  OR2 C2869 ( .A(n287), .B(n286), .Z(N790) );
  OR2 C2872 ( .A(N743), .B(N790), .Z(N7911) );
  OR2 C2874 ( .A(N7911), .B(N295), .Z(N792) );
  OR2 C2887 ( .A(N7911), .B(N740), .Z(N794) );
  OR2 C2900 ( .A(N7911), .B(N747), .Z(N796) );
  OR2 C2914 ( .A(N7911), .B(N750), .Z(N798) );
  OR2 C2927 ( .A(N7911), .B(N754), .Z(N800) );
  OR2 C2941 ( .A(N7911), .B(N757), .Z(N802) );
  OR2 C2955 ( .A(N7911), .B(N760), .Z(N804) );
  OR2 C2970 ( .A(N7911), .B(N764), .Z(N806) );
  OR2 C2983 ( .A(N7911), .B(N768), .Z(N808) );
  OR2 C2997 ( .A(N7911), .B(N7711), .Z(N8101) );
  OR2 C3011 ( .A(N7911), .B(N774), .Z(N8121) );
  OR2 C3025 ( .A(N767), .B(N763), .Z(N814) );
  OR2 C3026 ( .A(N7911), .B(N814), .Z(N815) );
  OR2 C3040 ( .A(N7911), .B(N779), .Z(N817) );
  OR2 C3054 ( .A(N786), .B(N739), .Z(N819) );
  OR2 C3055 ( .A(N7911), .B(N819), .Z(N820) );
  OR2 C3069 ( .A(N786), .B(N745), .Z(N822) );
  OR2 C3070 ( .A(N7911), .B(N822), .Z(N823) );
  AN2 C3072 ( .A(tx_8b_enc_in[7]), .B(tx_8b_enc_in[6]), .Z(N825) );
  AN2 C3073 ( .A(tx_8b_enc_in[5]), .B(tx_8b_enc_in[4]), .Z(N826) );
  AN2 C3074 ( .A(tx_8b_enc_in[3]), .B(tx_8b_enc_in[2]), .Z(N827) );
  AN2 C3075 ( .A(tx_8b_enc_in[1]), .B(tx_8b_enc_in[0]), .Z(N828) );
  AN2 C3076 ( .A(N825), .B(N826), .Z(N829) );
  AN2 C3077 ( .A(N827), .B(N828), .Z(N830) );
  AN2 C3078 ( .A(N829), .B(N830), .Z(N8311) );
  AN2 C5522 ( .A(n303), .B(n302), .Z(N842) );
  AN2 C5523 ( .A(n301), .B(n296), .Z(N843) );
  AN2 C5524 ( .A(N842), .B(N843), .Z(N844) );
  OR2 C5528 ( .A(N847), .B(N869), .Z(N845) );
  OR2 C5531 ( .A(encoder_sel[3]), .B(encoder_sel[2]), .Z(N847) );
  OR2 C5533 ( .A(N847), .B(N854), .Z(N848) );
  OR2 C5538 ( .A(N859), .B(N863), .Z(N850) );
  OR2 C5544 ( .A(N859), .B(N869), .Z(N852) );
  OR2 C5549 ( .A(n301), .B(encoder_sel[0]), .Z(N854) );
  OR2 C5550 ( .A(N859), .B(N854), .Z(N855) );
  OR2 C5555 ( .A(encoder_sel[3]), .B(n302), .Z(N859) );
  OR2 C5556 ( .A(n301), .B(n296), .Z(N860) );
  OR2 C5557 ( .A(N859), .B(N860), .Z(N8611) );
  OR2 C5561 ( .A(encoder_sel[1]), .B(encoder_sel[0]), .Z(N863) );
  OR2 C5562 ( .A(N868), .B(N863), .Z(N864) );
  OR2 C5566 ( .A(n303), .B(encoder_sel[2]), .Z(N868) );
  OR2 C5567 ( .A(encoder_sel[1]), .B(n296), .Z(N869) );
  OR2 C5568 ( .A(N868), .B(N869), .Z(N870) );
  OR2 C5721 ( .A(n165), .B(n175), .Z(N904) );
  OR2 C5739 ( .A(n34), .B(n154), .Z(N922) );
  OR2 C5885 ( .A(n157), .B(n168), .Z(N9911) );
  OR2 C6002 ( .A(n161), .B(n168), .Z(N1097) );
  OR2 C6022 ( .A(n161), .B(n157), .Z(N1116) );
  OR2 C6061 ( .A(n40), .B(n37), .Z(N1154) );
  OR2 C6086 ( .A(n294), .B(n292), .Z(N1177) );
  OR2 C6090 ( .A(n299), .B(n297), .Z(N1180) );
  IV I_04 ( .A(reset_tx), .Z(N213) );
  IV I_03 ( .A(reset_tx), .Z(N212) );
  AN2 C6 ( .A(N411), .B(N511), .Z(N611) );
  OR2 C8 ( .A(txd_sel[1]), .B(N511), .Z(N711) );
  OR2 C11 ( .A(N411), .B(txd_sel[0]), .Z(N911) );
  IV I_02 ( .A(txd_sel[1]), .Z(N411) );
  IV I_110 ( .A(txd_sel[0]), .Z(N511) );
  IV I_210 ( .A(N711), .Z(N811) );
  IV I_310 ( .A(N911), .Z(N1011) );
  IV I_01 ( .A(reset_tx), .Z(N210) );
  OR2 C128 ( .A(N20), .B(N25), .Z(N109) );
  OR2 C127 ( .A(N109), .B(N31), .Z(N110) );
  OR2 C126 ( .A(N110), .B(N36), .Z(N111) );
  OR2 C125 ( .A(N111), .B(N42), .Z(N112) );
  OR2 C124 ( .A(N112), .B(N49), .Z(N113) );
  AN2 C123 ( .A(N12), .B(N14), .Z(N106) );
  AN2 C122 ( .A(N106), .B(link_up_loc), .Z(N107) );
  AN2 C121 ( .A(N107), .B(N16), .Z(N108) );
  AN2 C120 ( .A(N108), .B(N113), .Z(assertion_shengyushen) );
  AN2 C119 ( .A(tx_er_d), .B(n14), .Z(txd_eq_crs_ext) );
  OR2 C118 ( .A(n4), .B(n5), .Z(N99) );
  OR2 C117 ( .A(N99), .B(n6), .Z(N100) );
  OR2 C116 ( .A(N100), .B(n7), .Z(N101) );
  OR2 C115 ( .A(N101), .B(n8), .Z(N102) );
  OR2 C114 ( .A(N102), .B(n9), .Z(N103) );
  OR2 C113 ( .A(N103), .B(n10), .Z(N104) );
  OR2 C112 ( .A(N104), .B(n1), .Z(N105) );
  OR2 C111 ( .A(N105), .B(n2), .Z(special_char) );
  OR2 C107 ( .A(n13), .B(N96), .Z(N97) );
  OR2 C106 ( .A(tx_enc_sel[1]), .B(N95), .Z(N96) );
  OR2 C105 ( .A(tx_enc_sel[2]), .B(n3), .Z(N95) );
  OR2 C101 ( .A(tx_enc_sel[0]), .B(N90), .Z(N91) );
  OR2 C100 ( .A(tx_enc_sel[1]), .B(N89), .Z(N90) );
  OR2 C99 ( .A(tx_enc_sel[2]), .B(n3), .Z(N89) );
  OR2 C96 ( .A(tx_enc_sel[0]), .B(N85), .Z(N86) );
  OR2 C95 ( .A(n12), .B(N84), .Z(N85) );
  OR2 C94 ( .A(n11), .B(tx_enc_sel[3]), .Z(N84) );
  OR2 C90 ( .A(n13), .B(N79), .Z(N80) );
  OR2 C89 ( .A(n12), .B(N78), .Z(N79) );
  OR2 C88 ( .A(n11), .B(tx_enc_sel[3]), .Z(N78) );
  OR2 C83 ( .A(n13), .B(N72), .Z(N73) );
  OR2 C82 ( .A(tx_enc_sel[1]), .B(N71), .Z(N72) );
  OR2 C81 ( .A(n11), .B(tx_enc_sel[3]), .Z(N71) );
  OR2 C77 ( .A(tx_enc_sel[0]), .B(N66), .Z(N67) );
  OR2 C76 ( .A(tx_enc_sel[1]), .B(N65), .Z(N66) );
  OR2 C75 ( .A(n11), .B(tx_enc_sel[3]), .Z(N65) );
  OR2 C72 ( .A(tx_enc_sel[0]), .B(N61), .Z(N62) );
  OR2 C71 ( .A(n12), .B(N60), .Z(N61) );
  OR2 C70 ( .A(tx_enc_sel[2]), .B(tx_enc_sel[3]), .Z(N60) );
  OR2 C67 ( .A(n13), .B(N56), .Z(N57) );
  OR2 C66 ( .A(tx_enc_sel[1]), .B(N55), .Z(N56) );
  OR2 C65 ( .A(tx_enc_sel[2]), .B(tx_enc_sel[3]), .Z(N55) );
  OR2 C62 ( .A(tx_enc_sel[0]), .B(N51), .Z(N52) );
  OR2 C61 ( .A(tx_enc_sel[1]), .B(N50), .Z(N51) );
  OR2 C60 ( .A(tx_enc_sel[2]), .B(tx_enc_sel[3]), .Z(N50) );
  IV I_22 ( .A(N48), .Z(N49) );
  OR2 C58 ( .A(N45), .B(N47), .Z(N48) );
  OR2 C57 ( .A(N44), .B(N46), .Z(N47) );
  OR2 C56 ( .A(N43), .B(tx_enc_ctrl_sel[3]), .Z(N46) );
  IV I_21 ( .A(tx_enc_ctrl_sel[0]), .Z(N45) );
  IV I_20 ( .A(tx_enc_ctrl_sel[1]), .Z(N44) );
  IV I_19 ( .A(tx_enc_ctrl_sel[2]), .Z(N43) );
  IV I_18 ( .A(N41), .Z(N42) );
  OR2 C51 ( .A(N38), .B(N40), .Z(N41) );
  OR2 C50 ( .A(tx_enc_ctrl_sel[1]), .B(N39), .Z(N40) );
  OR2 C49 ( .A(N37), .B(tx_enc_ctrl_sel[3]), .Z(N39) );
  IV I_17 ( .A(tx_enc_ctrl_sel[0]), .Z(N38) );
  IV I_16 ( .A(tx_enc_ctrl_sel[2]), .Z(N37) );
  IV I_15 ( .A(N35), .Z(N36) );
  OR2 C45 ( .A(tx_enc_ctrl_sel[0]), .B(N34), .Z(N35) );
  OR2 C44 ( .A(tx_enc_ctrl_sel[1]), .B(N33), .Z(N34) );
  OR2 C43 ( .A(N32), .B(tx_enc_ctrl_sel[3]), .Z(N33) );
  IV I_14 ( .A(tx_enc_ctrl_sel[2]), .Z(N32) );
  IV I_13 ( .A(N30), .Z(N31) );
  OR2 C40 ( .A(N27), .B(N29), .Z(N30) );
  OR2 C39 ( .A(N26), .B(N28), .Z(N29) );
  OR2 C38 ( .A(tx_enc_ctrl_sel[2]), .B(tx_enc_ctrl_sel[3]), .Z(N28) );
  IV I_12 ( .A(tx_enc_ctrl_sel[0]), .Z(N27) );
  IV I_11 ( .A(tx_enc_ctrl_sel[1]), .Z(N26) );
  IV I_10 ( .A(N24), .Z(N25) );
  OR2 C34 ( .A(tx_enc_ctrl_sel[0]), .B(N23), .Z(N24) );
  OR2 C33 ( .A(N21), .B(N22), .Z(N23) );
  OR2 C32 ( .A(tx_enc_ctrl_sel[2]), .B(tx_enc_ctrl_sel[3]), .Z(N22) );
  IV I_9 ( .A(tx_enc_ctrl_sel[1]), .Z(N21) );
  IV I_8 ( .A(N19), .Z(N20) );
  OR2 C29 ( .A(tx_enc_ctrl_sel[0]), .B(N18), .Z(N19) );
  OR2 C28 ( .A(tx_enc_ctrl_sel[1]), .B(N17), .Z(N18) );
  OR2 C27 ( .A(tx_enc_ctrl_sel[2]), .B(tx_enc_ctrl_sel[3]), .Z(N17) );
  IV I_7 ( .A(N15), .Z(N16) );
  OR2 C25 ( .A(jitter_study_pci[0]), .B(jitter_study_pci[1]), .Z(N15) );
  IV I_6 ( .A(N13), .Z(N14) );
  OR2 C23 ( .A(txd_sel[0]), .B(txd_sel[1]), .Z(N13) );
  IV I_5 ( .A(reset_tx), .Z(N12) );
  OR2 C20 ( .A(n15), .B(N9), .Z(N10) );
  OR2 C19 ( .A(n16), .B(N8), .Z(N9) );
  OR2 C18 ( .A(n17), .B(N7), .Z(N8) );
  OR2 C17 ( .A(n18), .B(N6), .Z(N7) );
  OR2 C16 ( .A(txd_d[4]), .B(N5), .Z(N6) );
  OR2 C15 ( .A(txd_d[5]), .B(N4), .Z(N5) );
  OR2 C14 ( .A(txd_d[6]), .B(txd_d[7]), .Z(N4) );
  FD1 qout_reg_0_ ( .D(n3399), .CP(txclk), .Q(txd_d[0]) );
  FD1 qout_reg_1_ ( .D(n3400), .CP(txclk), .Q(txd_d[1]) );
  FD1 qout_reg_2_ ( .D(n3401), .CP(txclk), .Q(txd_d[2]) );
  FD1 qout_reg_3_ ( .D(n3402), .CP(txclk), .Q(txd_d[3]) );
  FD1 qout_reg_4_ ( .D(n3403), .CP(txclk), .Q(txd_d[4]) );
  FD1 qout_reg_5_ ( .D(n3404), .CP(txclk), .Q(txd_d[5]) );
  FD1 qout_reg_6_ ( .D(n3405), .CP(txclk), .Q(txd_d[6]) );
  FD1 qout_reg_7_ ( .D(n3406), .CP(txclk), .Q(txd_d[7]) );
  FD1 qout_reg_0_1 ( .D(tx_8bdata_conf[0]), .CP(txclk), .Q(tx_8b_enc_in[0]) );
  FD1 qout_reg_1_1 ( .D(tx_8bdata_conf[1]), .CP(txclk), .Q(tx_8b_enc_in[1]) );
  FD1 qout_reg_2_1 ( .D(tx_8bdata_conf[2]), .CP(txclk), .Q(tx_8b_enc_in[2]) );
  FD1 qout_reg_3_1 ( .D(tx_8bdata_conf[3]), .CP(txclk), .Q(tx_8b_enc_in[3]) );
  FD1 qout_reg_4_1 ( .D(n3387), .CP(txclk), .Q(tx_8b_enc_in[4]) );
  FD1 qout_reg_5_1 ( .D(tx_8bdata_conf[5]), .CP(txclk), .Q(tx_8b_enc_in[5]) );
  FD1 qout_reg_6_1 ( .D(tx_8bdata_conf[6]), .CP(txclk), .Q(tx_8b_enc_in[6]) );
  FD1 qout_reg_7_1 ( .D(n3398), .CP(txclk), .Q(tx_8b_enc_in[7]) );
  FD1 qout_reg_0_2 ( .D(n3368), .CP(txclk), .Q(tx_en_d) );
  FD1 qout_reg_0_3 ( .D(n3367), .CP(txclk), .Q(tx_er_d) );
  FD1 qout_reg_0_4 ( .D(reset_tx), .CP(txclk), .Q(rst_reg) );
  FD1 qout_reg_0_8 ( .D(tx_enc_ctrl_sel[0]), .CP(txclk), .Q(
        tx_enc_ctrl_sel_reg[0]) );
  FD1 qout_reg_1_4 ( .D(tx_enc_ctrl_sel[1]), .CP(txclk), .Q(
        tx_enc_ctrl_sel_reg[1]) );
  FD1 qout_reg_2_4 ( .D(tx_enc_ctrl_sel[2]), .CP(txclk), .Q(
        tx_enc_ctrl_sel_reg[2]) );
  FD1 qout_reg_3_4 ( .D(tx_enc_ctrl_sel[3]), .CP(txclk), .Q(
        tx_enc_ctrl_sel_reg[3]) );
  FD1 qout_reg_0_9 ( .D(tx_enc_sel[0]), .CP(txclk), .Q(encoder_sel[0]) );
  FD1 qout_reg_1_5 ( .D(tx_enc_sel[1]), .CP(txclk), .Q(encoder_sel[1]) );
  FD1 qout_reg_2_5 ( .D(tx_enc_sel[2]), .CP(txclk), .Q(encoder_sel[2]) );
  FD1 qout_reg_3_5 ( .D(tx_enc_sel[3]), .CP(txclk), .Q(encoder_sel[3]) );
  FD1 qout_reg_0_10 ( .D(special_char), .CP(txclk), .Q(special_enc_in) );
  FD1 qout_reg_0_5 ( .D(n891), .CP(txclk), .Q(pos_disp_tx) );
  FD1 qout_reg_9_ ( .D(tx_10b_enc_out[9]), .CP(txclk), .Q(tx_10bdata_todiag[9]) );
  FD1 qout_reg_8_ ( .D(tx_10b_enc_out[8]), .CP(txclk), .Q(tx_10bdata_todiag[8]) );
  FD1 qout_reg_7_2 ( .D(tx_10b_enc_out[7]), .CP(txclk), .Q(
        tx_10bdata_todiag[7]) );
  FD1 qout_reg_6_2 ( .D(tx_10b_enc_out[6]), .CP(txclk), .Q(
        tx_10bdata_todiag[6]) );
  FD1 qout_reg_5_2 ( .D(tx_10b_enc_out[5]), .CP(txclk), .Q(
        tx_10bdata_todiag[5]) );
  FD1 qout_reg_4_2 ( .D(tx_10b_enc_out[4]), .CP(txclk), .Q(
        tx_10bdata_todiag[4]) );
  FD1 qout_reg_3_2 ( .D(tx_10b_enc_out[3]), .CP(txclk), .Q(
        tx_10bdata_todiag[3]) );
  FD1 qout_reg_2_2 ( .D(tx_10b_enc_out[2]), .CP(txclk), .Q(
        tx_10bdata_todiag[2]) );
  FD1 qout_reg_1_2 ( .D(tx_10b_enc_out[1]), .CP(txclk), .Q(
        tx_10bdata_todiag[1]) );
  FD1 qout_reg_0_6 ( .D(tx_10b_enc_out[0]), .CP(txclk), .Q(
        tx_10bdata_todiag[0]) );
  FD1 sync1_reg ( .D(jitter_study_pci[1]), .CP(txclk), .Q(sync1) );
  FD1 Q_reg ( .D(sync1), .CP(txclk), .Q(jitter_study_tx[1]) );
  FD1 sync1_reg1 ( .D(jitter_study_pci[0]), .CP(txclk), .Q(sync11) );
  FD1 Q_reg1 ( .D(sync11), .CP(txclk), .Q(jitter_study_tx[0]) );
  FD1 qout_reg_0_7 ( .D(n876), .CP(txclk), .Q(tx_10bdata[0]) );
  FD1 qout_reg_1_3 ( .D(n878), .CP(txclk), .Q(tx_10bdata[1]) );
  FD1 qout_reg_2_3 ( .D(n879), .CP(txclk), .Q(tx_10bdata[2]) );
  FD1 qout_reg_3_3 ( .D(tx_10bdata_predel[3]), .CP(txclk), .Q(tx_10bdata[3])
         );
  FD1 qout_reg_4_3 ( .D(tx_10bdata_predel[4]), .CP(txclk), .Q(tx_10bdata[4])
         );
  FD1 qout_reg_5_3 ( .D(tx_10bdata_predel[5]), .CP(txclk), .Q(tx_10bdata[5])
         );
  FD1 qout_reg_6_3 ( .D(tx_10bdata_predel[6]), .CP(txclk), .Q(tx_10bdata[6])
         );
  FD1 qout_reg_7_3 ( .D(tx_10bdata_predel[7]), .CP(txclk), .Q(tx_10bdata[7])
         );
  FD1 qout_reg_8_1 ( .D(n888), .CP(txclk), .Q(tx_10bdata[8]) );
  FD1 qout_reg_9_1 ( .D(n890), .CP(txclk), .Q(tx_10bdata[9]) );
  AN2 U870 ( .A(txd[7]), .B(N210), .Z(n3406) );
  AN2 U872 ( .A(txd[6]), .B(N210), .Z(n3405) );
  AN2 U874 ( .A(txd[5]), .B(N210), .Z(n3404) );
  AN2 U876 ( .A(txd[4]), .B(N210), .Z(n3403) );
  AN2 U878 ( .A(txd[3]), .B(N210), .Z(n3402) );
  AN2 U880 ( .A(txd[2]), .B(N210), .Z(n3401) );
  AN2 U882 ( .A(txd[1]), .B(N210), .Z(n3400) );
  AN2 U884 ( .A(txd[0]), .B(N210), .Z(n3399) );
  OR2 U885 ( .A(n3396), .B(n3397), .Z(n3398) );
  AN2 U886 ( .A(adver_reg[7]), .B(N811), .Z(n3397) );
  AN2 U887 ( .A(txd_d[7]), .B(N611), .Z(n3396) );
  OR2 U888 ( .A(n3395), .B(n3394), .Z(tx_8bdata_conf[6]) );
  OR2 U889 ( .A(n3392), .B(n3393), .Z(n3395) );
  AN2 U890 ( .A(ack), .B(N1011), .Z(n3394) );
  AN2 U891 ( .A(adver_reg[6]), .B(N811), .Z(n3393) );
  AN2 U892 ( .A(txd_d[6]), .B(N611), .Z(n3392) );
  OR2 U893 ( .A(n3391), .B(n3390), .Z(tx_8bdata_conf[5]) );
  OR2 U894 ( .A(n3388), .B(n3389), .Z(n3391) );
  AN2 U895 ( .A(adver_reg[12]), .B(N1011), .Z(n3390) );
  AN2 U896 ( .A(adver_reg[5]), .B(N811), .Z(n3389) );
  AN2 U897 ( .A(txd_d[5]), .B(N611), .Z(n3388) );
  OR2 U898 ( .A(n3385), .B(n3386), .Z(n3387) );
  AN2 U899 ( .A(adver_reg[4]), .B(N811), .Z(n3386) );
  AN2 U900 ( .A(txd_d[4]), .B(N611), .Z(n3385) );
  OR2 U901 ( .A(n3384), .B(n3383), .Z(tx_8bdata_conf[3]) );
  OR2 U902 ( .A(n3381), .B(n3382), .Z(n3384) );
  AN2 U903 ( .A(adver_reg[11]), .B(N1011), .Z(n3383) );
  AN2 U904 ( .A(adver_reg[3]), .B(N811), .Z(n3382) );
  AN2 U905 ( .A(txd_d[3]), .B(N611), .Z(n3381) );
  OR2 U906 ( .A(n3380), .B(n3379), .Z(tx_8bdata_conf[2]) );
  OR2 U907 ( .A(n3377), .B(n3378), .Z(n3380) );
  AN2 U908 ( .A(adver_reg[10]), .B(N1011), .Z(n3379) );
  AN2 U909 ( .A(adver_reg[2]), .B(N811), .Z(n3378) );
  AN2 U910 ( .A(txd_d[2]), .B(N611), .Z(n3377) );
  OR2 U911 ( .A(n3376), .B(n3375), .Z(tx_8bdata_conf[1]) );
  OR2 U912 ( .A(n3373), .B(n3374), .Z(n3376) );
  AN2 U913 ( .A(adver_reg[9]), .B(N1011), .Z(n3375) );
  AN2 U914 ( .A(adver_reg[1]), .B(N811), .Z(n3374) );
  AN2 U915 ( .A(txd_d[1]), .B(N611), .Z(n3373) );
  OR2 U916 ( .A(n3372), .B(n3371), .Z(tx_8bdata_conf[0]) );
  OR2 U917 ( .A(n3369), .B(n3370), .Z(n3372) );
  AN2 U918 ( .A(adver_reg[8]), .B(N1011), .Z(n3371) );
  AN2 U919 ( .A(adver_reg[0]), .B(N811), .Z(n3370) );
  AN2 U920 ( .A(txd_d[0]), .B(N611), .Z(n3369) );
  AN2 U922 ( .A(tx_en), .B(N212), .Z(n3368) );
  AN2 U924 ( .A(tx_er), .B(N213), .Z(n3367) );
  OR2 U925 ( .A(n3365), .B(n3366), .Z(tx_10b_enc_out[9]) );
  AN2 U926 ( .A(n3346), .B(special_enc_in), .Z(n3366) );
  AN2 U927 ( .A(N8411), .B(n304), .Z(n3365) );
  OR2 U928 ( .A(n3363), .B(n3364), .Z(tx_10b_enc_out[8]) );
  AN2 U929 ( .A(N889), .B(special_enc_in), .Z(n3364) );
  AN2 U930 ( .A(N840), .B(n304), .Z(n3363) );
  OR2 U931 ( .A(n3361), .B(n3362), .Z(tx_10b_enc_out[7]) );
  AN2 U932 ( .A(n3332), .B(special_enc_in), .Z(n3362) );
  AN2 U933 ( .A(N839), .B(n304), .Z(n3361) );
  OR2 U934 ( .A(n3359), .B(n3360), .Z(tx_10b_enc_out[6]) );
  AN2 U935 ( .A(N887), .B(special_enc_in), .Z(n3360) );
  AN2 U936 ( .A(N838), .B(n304), .Z(n3359) );
  OR2 U937 ( .A(n3357), .B(n3358), .Z(tx_10b_enc_out[5]) );
  AN2 U938 ( .A(N886), .B(special_enc_in), .Z(n3358) );
  AN2 U939 ( .A(N837), .B(n304), .Z(n3357) );
  OR2 U940 ( .A(n3355), .B(n3356), .Z(tx_10b_enc_out[4]) );
  AN2 U941 ( .A(N885), .B(special_enc_in), .Z(n3356) );
  AN2 U942 ( .A(N836), .B(n304), .Z(n3355) );
  OR2 U943 ( .A(n3353), .B(n3354), .Z(tx_10b_enc_out[3]) );
  AN2 U944 ( .A(N884), .B(special_enc_in), .Z(n3354) );
  AN2 U945 ( .A(N835), .B(n304), .Z(n3353) );
  OR2 U946 ( .A(n3351), .B(n3352), .Z(tx_10b_enc_out[2]) );
  AN2 U947 ( .A(N883), .B(special_enc_in), .Z(n3352) );
  AN2 U948 ( .A(N834), .B(n304), .Z(n3351) );
  OR2 U949 ( .A(n3349), .B(n3350), .Z(tx_10b_enc_out[1]) );
  AN2 U950 ( .A(N882), .B(special_enc_in), .Z(n3350) );
  AN2 U951 ( .A(N833), .B(n304), .Z(n3349) );
  OR2 U952 ( .A(n3347), .B(n3348), .Z(tx_10b_enc_out[0]) );
  AN2 U953 ( .A(N8811), .B(special_enc_in), .Z(n3348) );
  AN2 U954 ( .A(N832), .B(n304), .Z(n3347) );
  OR2 U955 ( .A(n3344), .B(n3345), .Z(n3346) );
  OR2 U956 ( .A(n3342), .B(n3343), .Z(n3345) );
  OR2 U957 ( .A(n3340), .B(n3341), .Z(n3344) );
  OR2 U958 ( .A(n3338), .B(n3339), .Z(n3343) );
  OR2 U959 ( .A(n3337), .B(N1180), .Z(n3342) );
  OR2 U960 ( .A(n3335), .B(n3336), .Z(n3341) );
  OR2 U961 ( .A(n3333), .B(n3334), .Z(n3340) );
  AN2 U962 ( .A(n291), .B(n292), .Z(n3339) );
  AN2 U963 ( .A(pos_disp_tx), .B(n295), .Z(n3338) );
  AN2 U964 ( .A(n291), .B(n293), .Z(n3337) );
  AN2 U965 ( .A(n291), .B(n298), .Z(n3336) );
  AN2 U966 ( .A(n291), .B(n300), .Z(n3335) );
  AN2 U967 ( .A(pos_disp_tx), .B(n294), .Z(n3334) );
  AN2 U968 ( .A(pos_disp_tx), .B(N844), .Z(n3333) );
  OR2 U969 ( .A(n3330), .B(n3331), .Z(n3332) );
  OR2 U970 ( .A(n3328), .B(n3329), .Z(n3331) );
  OR2 U971 ( .A(n3326), .B(n3327), .Z(n3330) );
  OR2 U972 ( .A(n3324), .B(n3325), .Z(n3329) );
  OR2 U973 ( .A(n3323), .B(N1180), .Z(n3328) );
  OR2 U974 ( .A(n3321), .B(n3322), .Z(n3327) );
  OR2 U975 ( .A(n3319), .B(n3320), .Z(n3326) );
  AN2 U976 ( .A(n291), .B(n292), .Z(n3325) );
  AN2 U977 ( .A(n291), .B(n295), .Z(n3324) );
  AN2 U978 ( .A(n291), .B(n293), .Z(n3323) );
  AN2 U979 ( .A(n291), .B(n298), .Z(n3322) );
  AN2 U980 ( .A(pos_disp_tx), .B(n300), .Z(n3321) );
  AN2 U981 ( .A(n291), .B(n294), .Z(n3320) );
  AN2 U982 ( .A(n291), .B(N844), .Z(n3319) );
  OR2 U983 ( .A(n3317), .B(n3318), .Z(N889) );
  OR2 U984 ( .A(n3311), .B(n3316), .Z(n3318) );
  OR2 U985 ( .A(n3314), .B(n3315), .Z(n3317) );
  OR2 U986 ( .A(n3312), .B(n3313), .Z(n3316) );
  OR2 U987 ( .A(n3309), .B(n3310), .Z(n3315) );
  OR2 U988 ( .A(n3307), .B(n3308), .Z(n3314) );
  AN2 U989 ( .A(pos_disp_tx), .B(n292), .Z(n3313) );
  AN2 U990 ( .A(n291), .B(n295), .Z(n3312) );
  AN2 U991 ( .A(n291), .B(n293), .Z(n3311) );
  AN2 U992 ( .A(pos_disp_tx), .B(n298), .Z(n3310) );
  AN2 U993 ( .A(n291), .B(n300), .Z(n3309) );
  AN2 U994 ( .A(n291), .B(n294), .Z(n3308) );
  AN2 U995 ( .A(pos_disp_tx), .B(N844), .Z(n3307) );
  OR2 U996 ( .A(n3305), .B(n3306), .Z(N887) );
  OR2 U997 ( .A(n3299), .B(n3304), .Z(n3306) );
  OR2 U998 ( .A(n3302), .B(n3303), .Z(n3305) );
  OR2 U999 ( .A(n3300), .B(n3301), .Z(n3304) );
  OR2 U1000 ( .A(n3297), .B(n3298), .Z(n3303) );
  OR2 U1001 ( .A(n3295), .B(n3296), .Z(n3302) );
  AN2 U1002 ( .A(n291), .B(n292), .Z(n3301) );
  AN2 U1003 ( .A(n291), .B(n295), .Z(n3300) );
  AN2 U1004 ( .A(pos_disp_tx), .B(n293), .Z(n3299) );
  AN2 U1005 ( .A(n291), .B(n298), .Z(n3298) );
  AN2 U1006 ( .A(n291), .B(n300), .Z(n3297) );
  AN2 U1007 ( .A(pos_disp_tx), .B(n294), .Z(n3296) );
  AN2 U1008 ( .A(n291), .B(N844), .Z(n3295) );
  OR2 U1009 ( .A(n3294), .B(n3288), .Z(N886) );
  OR2 U1010 ( .A(n3292), .B(n3293), .Z(n3294) );
  OR2 U1011 ( .A(n3286), .B(n3291), .Z(n3293) );
  OR2 U1012 ( .A(n3289), .B(n3290), .Z(n3292) );
  OR2 U1013 ( .A(n3287), .B(n297), .Z(n3291) );
  OR2 U1014 ( .A(n3284), .B(n3285), .Z(n3290) );
  OR2 U1015 ( .A(n3282), .B(n3283), .Z(n3289) );
  AN2 U1016 ( .A(pos_disp_tx), .B(n292), .Z(n3288) );
  AN2 U1017 ( .A(n291), .B(n295), .Z(n3287) );
  AN2 U1018 ( .A(n291), .B(n293), .Z(n3286) );
  AN2 U1019 ( .A(n291), .B(n298), .Z(n3285) );
  AN2 U1020 ( .A(n291), .B(n300), .Z(n3284) );
  AN2 U1021 ( .A(n291), .B(n294), .Z(n3283) );
  AN2 U1022 ( .A(n291), .B(N844), .Z(n3282) );
  OR2 U1023 ( .A(n3281), .B(n3275), .Z(N885) );
  OR2 U1024 ( .A(n3279), .B(n3280), .Z(n3281) );
  OR2 U1025 ( .A(n3278), .B(n3274), .Z(n3280) );
  OR2 U1026 ( .A(n3276), .B(n3277), .Z(n3279) );
  OR2 U1027 ( .A(n3273), .B(n299), .Z(n3278) );
  OR2 U1028 ( .A(n3271), .B(n3272), .Z(n3277) );
  OR2 U1029 ( .A(n3269), .B(n3270), .Z(n3276) );
  AN2 U1030 ( .A(n291), .B(n292), .Z(n3275) );
  AN2 U1031 ( .A(pos_disp_tx), .B(n295), .Z(n3274) );
  AN2 U1032 ( .A(pos_disp_tx), .B(n293), .Z(n3273) );
  AN2 U1033 ( .A(pos_disp_tx), .B(n298), .Z(n3272) );
  AN2 U1034 ( .A(pos_disp_tx), .B(n300), .Z(n3271) );
  AN2 U1035 ( .A(n291), .B(n294), .Z(n3270) );
  AN2 U1036 ( .A(n291), .B(N844), .Z(n3269) );
  OR2 U1037 ( .A(n3267), .B(n3268), .Z(N884) );
  OR2 U1038 ( .A(n3266), .B(n297), .Z(n3268) );
  OR2 U1039 ( .A(n3260), .B(n3265), .Z(n3267) );
  OR2 U1040 ( .A(n3263), .B(n3264), .Z(n3266) );
  OR2 U1041 ( .A(n3261), .B(n3262), .Z(n3265) );
  AN2 U1042 ( .A(n291), .B(n295), .Z(n3264) );
  AN2 U1043 ( .A(n291), .B(n293), .Z(n3263) );
  AN2 U1044 ( .A(n291), .B(n298), .Z(n3262) );
  AN2 U1045 ( .A(n291), .B(n300), .Z(n3261) );
  AN2 U1046 ( .A(n291), .B(N844), .Z(n3260) );
  OR2 U1047 ( .A(n3259), .B(n3258), .Z(N883) );
  OR2 U1048 ( .A(n3256), .B(n3257), .Z(n3259) );
  OR2 U1049 ( .A(n3254), .B(n3255), .Z(n3258) );
  OR2 U1050 ( .A(n3252), .B(n3253), .Z(n3257) );
  OR2 U1051 ( .A(n3251), .B(N11811), .Z(n3256) );
  AN2 U1052 ( .A(pos_disp_tx), .B(n295), .Z(n3255) );
  AN2 U1053 ( .A(pos_disp_tx), .B(n293), .Z(n3254) );
  AN2 U1054 ( .A(pos_disp_tx), .B(n298), .Z(n3253) );
  AN2 U1055 ( .A(pos_disp_tx), .B(n300), .Z(n3252) );
  AN2 U1056 ( .A(pos_disp_tx), .B(N844), .Z(n3251) );
  OR2 U1057 ( .A(n3249), .B(n3250), .Z(N882) );
  OR2 U1058 ( .A(n3248), .B(n3246), .Z(n3250) );
  OR2 U1059 ( .A(n3242), .B(n3247), .Z(n3249) );
  OR2 U1060 ( .A(n3245), .B(N1180), .Z(n3248) );
  OR2 U1061 ( .A(n3243), .B(n3244), .Z(n3247) );
  AN2 U1062 ( .A(pos_disp_tx), .B(n295), .Z(n3246) );
  AN2 U1063 ( .A(pos_disp_tx), .B(n293), .Z(n3245) );
  AN2 U1064 ( .A(pos_disp_tx), .B(n298), .Z(n3244) );
  AN2 U1065 ( .A(pos_disp_tx), .B(n300), .Z(n3243) );
  AN2 U1066 ( .A(n291), .B(N844), .Z(n3242) );
  OR2 U1067 ( .A(n3240), .B(n3241), .Z(N8811) );
  OR2 U1068 ( .A(n3236), .B(n3237), .Z(n3241) );
  OR2 U1069 ( .A(n3238), .B(n3239), .Z(n3240) );
  OR2 U1070 ( .A(n3234), .B(n3235), .Z(n3239) );
  OR2 U1071 ( .A(n3233), .B(N1177), .Z(n3238) );
  AN2 U1072 ( .A(pos_disp_tx), .B(n295), .Z(n3237) );
  AN2 U1073 ( .A(pos_disp_tx), .B(n293), .Z(n3236) );
  AN2 U1074 ( .A(pos_disp_tx), .B(n298), .Z(n3235) );
  AN2 U1075 ( .A(pos_disp_tx), .B(n300), .Z(n3234) );
  AN2 U1076 ( .A(pos_disp_tx), .B(N844), .Z(n3233) );
  OR2 U1077 ( .A(n3231), .B(n3232), .Z(N8411) );
  OR2 U1078 ( .A(n3229), .B(n3230), .Z(n3232) );
  OR2 U1079 ( .A(n3227), .B(n3228), .Z(n3231) );
  OR2 U1080 ( .A(n3226), .B(n3177), .Z(n3230) );
  OR2 U1081 ( .A(n3224), .B(n3225), .Z(n3229) );
  OR2 U1082 ( .A(n3222), .B(n3223), .Z(n3228) );
  OR2 U1083 ( .A(n3220), .B(n3221), .Z(n3227) );
  OR2 U1084 ( .A(n3218), .B(n3219), .Z(n3226) );
  OR2 U1085 ( .A(n3216), .B(n3217), .Z(n3225) );
  OR2 U1086 ( .A(n3214), .B(n3215), .Z(n3224) );
  OR2 U1087 ( .A(n3212), .B(n3213), .Z(n3223) );
  OR2 U1088 ( .A(n3210), .B(n3211), .Z(n3222) );
  OR2 U1089 ( .A(n3208), .B(n3209), .Z(n3221) );
  OR2 U1090 ( .A(n3206), .B(n3207), .Z(n3220) );
  OR2 U1091 ( .A(n3204), .B(n3205), .Z(n3219) );
  OR2 U1092 ( .A(n3202), .B(n3203), .Z(n3218) );
  OR2 U1093 ( .A(n3200), .B(n3201), .Z(n3217) );
  OR2 U1094 ( .A(n3198), .B(n3199), .Z(n3216) );
  OR2 U1095 ( .A(n3196), .B(n3197), .Z(n3215) );
  OR2 U1096 ( .A(n3194), .B(n3195), .Z(n3214) );
  OR2 U1097 ( .A(n3192), .B(n3193), .Z(n3213) );
  OR2 U1098 ( .A(n3190), .B(n3191), .Z(n3212) );
  OR2 U1099 ( .A(n3188), .B(n3189), .Z(n3211) );
  OR2 U1100 ( .A(n3186), .B(n3187), .Z(n3210) );
  OR2 U1101 ( .A(n3184), .B(n3185), .Z(n3209) );
  OR2 U1102 ( .A(n3182), .B(n3183), .Z(n3208) );
  OR2 U1103 ( .A(n3180), .B(n3181), .Z(n3207) );
  OR2 U1104 ( .A(n3178), .B(n3179), .Z(n3206) );
  OR2 U1105 ( .A(n3175), .B(n3176), .Z(n3205) );
  OR2 U1106 ( .A(n3173), .B(n3174), .Z(n3204) );
  OR2 U1107 ( .A(n3171), .B(n3172), .Z(n3203) );
  OR2 U1108 ( .A(n3169), .B(n3170), .Z(n3202) );
  OR2 U1109 ( .A(n3167), .B(n3168), .Z(n3201) );
  OR2 U1110 ( .A(n3165), .B(n3166), .Z(n3200) );
  OR2 U1111 ( .A(n3163), .B(n3164), .Z(n3199) );
  OR2 U1112 ( .A(n3161), .B(n3162), .Z(n3198) );
  OR2 U1113 ( .A(n3159), .B(n3160), .Z(n3197) );
  OR2 U1114 ( .A(n3157), .B(n3158), .Z(n3196) );
  OR2 U1115 ( .A(n3155), .B(n3156), .Z(n3195) );
  OR2 U1116 ( .A(n3153), .B(n3154), .Z(n3194) );
  OR2 U1117 ( .A(n3151), .B(n3152), .Z(n3193) );
  OR2 U1118 ( .A(n3149), .B(n3150), .Z(n3192) );
  OR2 U1119 ( .A(n3147), .B(n3148), .Z(n3191) );
  OR2 U1120 ( .A(n3145), .B(n3146), .Z(n3190) );
  OR2 U1121 ( .A(n3143), .B(n3144), .Z(n3189) );
  OR2 U1122 ( .A(n3141), .B(n3142), .Z(n3188) );
  OR2 U1123 ( .A(n3139), .B(n3140), .Z(n3187) );
  OR2 U1124 ( .A(n3137), .B(n3138), .Z(n3186) );
  OR2 U1125 ( .A(n3135), .B(n3136), .Z(n3185) );
  OR2 U1126 ( .A(n3133), .B(n3134), .Z(n3184) );
  OR2 U1127 ( .A(n3131), .B(n3132), .Z(n3183) );
  OR2 U1128 ( .A(n3129), .B(n3130), .Z(n3182) );
  OR2 U1129 ( .A(n3127), .B(n3128), .Z(n3181) );
  OR2 U1130 ( .A(n3125), .B(n3126), .Z(n3180) );
  OR2 U1131 ( .A(n3013), .B(n3124), .Z(n3179) );
  OR2 U1132 ( .A(n3122), .B(n3123), .Z(n3178) );
  OR2 U1133 ( .A(n3120), .B(n3121), .Z(n3177) );
  OR2 U1134 ( .A(n3118), .B(n3119), .Z(n3176) );
  OR2 U1135 ( .A(n3116), .B(n3117), .Z(n3175) );
  OR2 U1136 ( .A(n3114), .B(n3115), .Z(n3174) );
  OR2 U1137 ( .A(n3112), .B(n3113), .Z(n3173) );
  OR2 U1138 ( .A(n3110), .B(n3111), .Z(n3172) );
  OR2 U1139 ( .A(n3108), .B(n3109), .Z(n3171) );
  OR2 U1140 ( .A(n3106), .B(n3107), .Z(n3170) );
  OR2 U1141 ( .A(n3104), .B(n3105), .Z(n3169) );
  OR2 U1142 ( .A(n3102), .B(n3103), .Z(n3168) );
  OR2 U1143 ( .A(n3100), .B(n3101), .Z(n3167) );
  OR2 U1144 ( .A(n3098), .B(n3099), .Z(n3166) );
  OR2 U1145 ( .A(n3096), .B(n3097), .Z(n3165) );
  OR2 U1146 ( .A(n3094), .B(n3095), .Z(n3164) );
  OR2 U1147 ( .A(n3092), .B(n3093), .Z(n3163) );
  OR2 U1148 ( .A(n3090), .B(n3091), .Z(n3162) );
  OR2 U1149 ( .A(n3088), .B(n3089), .Z(n3161) );
  OR2 U1150 ( .A(n3086), .B(n3087), .Z(n3160) );
  OR2 U1151 ( .A(n3084), .B(n3085), .Z(n3159) );
  OR2 U1152 ( .A(n3082), .B(n3083), .Z(n3158) );
  OR2 U1153 ( .A(n3080), .B(n3081), .Z(n3157) );
  OR2 U1154 ( .A(n3078), .B(n3079), .Z(n3156) );
  OR2 U1155 ( .A(n3076), .B(n3077), .Z(n3155) );
  OR2 U1156 ( .A(n3074), .B(n3075), .Z(n3154) );
  OR2 U1157 ( .A(n3072), .B(n3073), .Z(n3153) );
  OR2 U1158 ( .A(n3070), .B(n3071), .Z(n3152) );
  OR2 U1159 ( .A(n3068), .B(n3069), .Z(n3151) );
  OR2 U1160 ( .A(n3066), .B(n3067), .Z(n3150) );
  OR2 U1161 ( .A(n3064), .B(n3065), .Z(n3149) );
  OR2 U1162 ( .A(n3062), .B(n3063), .Z(n3148) );
  OR2 U1163 ( .A(n3060), .B(n3061), .Z(n3147) );
  OR2 U1164 ( .A(n3058), .B(n3059), .Z(n3146) );
  OR2 U1165 ( .A(n3056), .B(n3057), .Z(n3145) );
  OR2 U1166 ( .A(n3054), .B(n3055), .Z(n3144) );
  OR2 U1167 ( .A(n3052), .B(n3053), .Z(n3143) );
  OR2 U1168 ( .A(n3050), .B(n3051), .Z(n3142) );
  OR2 U1169 ( .A(n3048), .B(n3049), .Z(n3141) );
  OR2 U1170 ( .A(n3046), .B(n3047), .Z(n3140) );
  OR2 U1171 ( .A(n3044), .B(n3045), .Z(n3139) );
  OR2 U1172 ( .A(n3042), .B(n3043), .Z(n3138) );
  OR2 U1173 ( .A(n3040), .B(n3041), .Z(n3137) );
  OR2 U1174 ( .A(n3038), .B(n3039), .Z(n3136) );
  OR2 U1175 ( .A(n3036), .B(n3037), .Z(n3135) );
  OR2 U1176 ( .A(n3034), .B(n3035), .Z(n3134) );
  OR2 U1177 ( .A(n3032), .B(n3033), .Z(n3133) );
  OR2 U1178 ( .A(n3030), .B(n3031), .Z(n3132) );
  OR2 U1179 ( .A(n3028), .B(n3029), .Z(n3131) );
  OR2 U1180 ( .A(n3026), .B(n3027), .Z(n3130) );
  OR2 U1181 ( .A(n3024), .B(n3025), .Z(n3129) );
  OR2 U1182 ( .A(n3022), .B(n3023), .Z(n3128) );
  OR2 U1183 ( .A(n3020), .B(n3021), .Z(n3127) );
  OR2 U1184 ( .A(n3018), .B(n3019), .Z(n3126) );
  OR2 U1185 ( .A(n3016), .B(n3017), .Z(n3125) );
  OR2 U1186 ( .A(n3014), .B(n3015), .Z(n3124) );
  OR2 U1187 ( .A(n3012), .B(N1158), .Z(n3123) );
  OR2 U1188 ( .A(n3010), .B(n3011), .Z(n3122) );
  AN2 U1189 ( .A(n291), .B(N8311), .Z(n3121) );
  AN2 U1190 ( .A(pos_disp_tx), .B(n153), .Z(n3120) );
  AN2 U1191 ( .A(n291), .B(n33), .Z(n3119) );
  AN2 U1192 ( .A(n291), .B(n19), .Z(n3118) );
  AN2 U1193 ( .A(n291), .B(n172), .Z(n3117) );
  AN2 U1194 ( .A(n291), .B(n26), .Z(n3116) );
  AN2 U1195 ( .A(pos_disp_tx), .B(n178), .Z(n3115) );
  AN2 U1196 ( .A(pos_disp_tx), .B(n23), .Z(n3114) );
  AN2 U1197 ( .A(n291), .B(n173), .Z(n3113) );
  AN2 U1198 ( .A(n291), .B(n27), .Z(n3112) );
  AN2 U1199 ( .A(n291), .B(n176), .Z(n3111) );
  AN2 U1200 ( .A(n291), .B(n166), .Z(n3110) );
  AN2 U1201 ( .A(pos_disp_tx), .B(n44), .Z(n3109) );
  AN2 U1202 ( .A(n291), .B(n179), .Z(n3108) );
  AN2 U1203 ( .A(n291), .B(n24), .Z(n3107) );
  AN2 U1204 ( .A(pos_disp_tx), .B(n155), .Z(n3106) );
  AN2 U1205 ( .A(n291), .B(n35), .Z(n3105) );
  AN2 U1206 ( .A(n291), .B(n21), .Z(n3104) );
  AN2 U1207 ( .A(n291), .B(n174), .Z(n3103) );
  AN2 U1208 ( .A(n291), .B(n28), .Z(n3102) );
  AN2 U1209 ( .A(pos_disp_tx), .B(n180), .Z(n3101) );
  AN2 U1210 ( .A(pos_disp_tx), .B(n25), .Z(n3100) );
  AN2 U1211 ( .A(n291), .B(n205), .Z(n3099) );
  AN2 U1212 ( .A(n291), .B(n29), .Z(n3098) );
  AN2 U1213 ( .A(n291), .B(n218), .Z(n3097) );
  AN2 U1214 ( .A(n291), .B(n267), .Z(n3096) );
  AN2 U1215 ( .A(pos_disp_tx), .B(n133), .Z(n3095) );
  AN2 U1216 ( .A(n291), .B(n181), .Z(n3094) );
  AN2 U1217 ( .A(n291), .B(n60), .Z(n3093) );
  AN2 U1218 ( .A(pos_disp_tx), .B(n231), .Z(n3092) );
  AN2 U1219 ( .A(n291), .B(n97), .Z(n3091) );
  AN2 U1220 ( .A(n291), .B(n48), .Z(n3090) );
  AN2 U1221 ( .A(n291), .B(n206), .Z(n3089) );
  AN2 U1222 ( .A(n291), .B(n72), .Z(n3088) );
  AN2 U1223 ( .A(pos_disp_tx), .B(n182), .Z(n3087) );
  AN2 U1224 ( .A(pos_disp_tx), .B(n61), .Z(n3086) );
  AN2 U1225 ( .A(n291), .B(n207), .Z(n3085) );
  AN2 U1226 ( .A(n291), .B(n73), .Z(n3084) );
  AN2 U1227 ( .A(n291), .B(n220), .Z(n3083) );
  AN2 U1228 ( .A(n291), .B(n269), .Z(n3082) );
  AN2 U1229 ( .A(pos_disp_tx), .B(n135), .Z(n3081) );
  AN2 U1230 ( .A(n291), .B(n183), .Z(n3080) );
  AN2 U1231 ( .A(n291), .B(n62), .Z(n3079) );
  AN2 U1232 ( .A(pos_disp_tx), .B(n233), .Z(n3078) );
  AN2 U1233 ( .A(n291), .B(n99), .Z(n3077) );
  AN2 U1234 ( .A(n291), .B(n50), .Z(n3076) );
  AN2 U1235 ( .A(n291), .B(n208), .Z(n3075) );
  AN2 U1236 ( .A(n291), .B(n74), .Z(n3074) );
  AN2 U1237 ( .A(pos_disp_tx), .B(n184), .Z(n3073) );
  AN2 U1238 ( .A(pos_disp_tx), .B(n63), .Z(n3072) );
  AN2 U1239 ( .A(n291), .B(n209), .Z(n3071) );
  AN2 U1240 ( .A(n291), .B(n75), .Z(n3070) );
  AN2 U1241 ( .A(n291), .B(n222), .Z(n3069) );
  AN2 U1242 ( .A(n291), .B(n271), .Z(n3068) );
  AN2 U1243 ( .A(pos_disp_tx), .B(n137), .Z(n3067) );
  AN2 U1244 ( .A(n291), .B(n185), .Z(n3066) );
  AN2 U1245 ( .A(n291), .B(n64), .Z(n3065) );
  AN2 U1246 ( .A(pos_disp_tx), .B(n235), .Z(n3064) );
  AN2 U1247 ( .A(n291), .B(n101), .Z(n3063) );
  AN2 U1248 ( .A(n291), .B(n52), .Z(n3062) );
  AN2 U1249 ( .A(n291), .B(n210), .Z(n3061) );
  AN2 U1250 ( .A(n291), .B(n76), .Z(n3060) );
  AN2 U1251 ( .A(pos_disp_tx), .B(n186), .Z(n3059) );
  AN2 U1252 ( .A(pos_disp_tx), .B(n65), .Z(n3058) );
  AN2 U1253 ( .A(n291), .B(n211), .Z(n3057) );
  AN2 U1254 ( .A(n291), .B(n77), .Z(n3056) );
  AN2 U1255 ( .A(n291), .B(n224), .Z(n3055) );
  AN2 U1256 ( .A(n291), .B(n273), .Z(n3054) );
  AN2 U1257 ( .A(pos_disp_tx), .B(n139), .Z(n3053) );
  AN2 U1258 ( .A(n291), .B(n187), .Z(n3052) );
  AN2 U1259 ( .A(n291), .B(n66), .Z(n3051) );
  AN2 U1260 ( .A(pos_disp_tx), .B(n237), .Z(n3050) );
  AN2 U1261 ( .A(n291), .B(n103), .Z(n3049) );
  AN2 U1262 ( .A(n291), .B(n54), .Z(n3048) );
  AN2 U1263 ( .A(n291), .B(n212), .Z(n3047) );
  AN2 U1264 ( .A(n291), .B(n78), .Z(n3046) );
  AN2 U1265 ( .A(pos_disp_tx), .B(n188), .Z(n3045) );
  AN2 U1266 ( .A(pos_disp_tx), .B(n67), .Z(n3044) );
  AN2 U1267 ( .A(n291), .B(n213), .Z(n3043) );
  AN2 U1268 ( .A(n291), .B(n79), .Z(n3042) );
  AN2 U1269 ( .A(n291), .B(n226), .Z(n3041) );
  AN2 U1270 ( .A(n291), .B(n275), .Z(n3040) );
  AN2 U1271 ( .A(pos_disp_tx), .B(n141), .Z(n3039) );
  AN2 U1272 ( .A(n291), .B(n189), .Z(n3038) );
  AN2 U1273 ( .A(n291), .B(n68), .Z(n3037) );
  AN2 U1274 ( .A(pos_disp_tx), .B(n239), .Z(n3036) );
  AN2 U1275 ( .A(n291), .B(n105), .Z(n3035) );
  AN2 U1276 ( .A(n291), .B(n56), .Z(n3034) );
  AN2 U1277 ( .A(n291), .B(n214), .Z(n3033) );
  AN2 U1278 ( .A(n291), .B(n80), .Z(n3032) );
  AN2 U1279 ( .A(pos_disp_tx), .B(n190), .Z(n3031) );
  AN2 U1280 ( .A(pos_disp_tx), .B(n69), .Z(n3030) );
  AN2 U1281 ( .A(n291), .B(n215), .Z(n3029) );
  AN2 U1282 ( .A(n291), .B(n81), .Z(n3028) );
  AN2 U1283 ( .A(n291), .B(n228), .Z(n3027) );
  AN2 U1284 ( .A(n291), .B(n277), .Z(n3026) );
  AN2 U1285 ( .A(pos_disp_tx), .B(n143), .Z(n3025) );
  AN2 U1286 ( .A(n291), .B(n191), .Z(n3024) );
  AN2 U1287 ( .A(n291), .B(n70), .Z(n3023) );
  AN2 U1288 ( .A(pos_disp_tx), .B(n241), .Z(n3022) );
  AN2 U1289 ( .A(n291), .B(n107), .Z(n3021) );
  AN2 U1290 ( .A(n291), .B(n58), .Z(n3020) );
  AN2 U1291 ( .A(n291), .B(n216), .Z(n3019) );
  AN2 U1292 ( .A(n291), .B(n82), .Z(n3018) );
  AN2 U1293 ( .A(pos_disp_tx), .B(n192), .Z(n3017) );
  AN2 U1294 ( .A(pos_disp_tx), .B(n71), .Z(n3016) );
  AN2 U1295 ( .A(n291), .B(n217), .Z(n3015) );
  AN2 U1296 ( .A(n291), .B(n83), .Z(n3014) );
  AN2 U1297 ( .A(n291), .B(n230), .Z(n3013) );
  AN2 U1298 ( .A(n291), .B(n279), .Z(n3012) );
  AN2 U1299 ( .A(pos_disp_tx), .B(n145), .Z(n3011) );
  AN2 U1300 ( .A(n291), .B(N239), .Z(n3010) );
  OR2 U1301 ( .A(n3008), .B(n3009), .Z(N840) );
  OR2 U1302 ( .A(n3006), .B(n3007), .Z(n3009) );
  OR2 U1303 ( .A(n3004), .B(n3005), .Z(n3008) );
  OR2 U1304 ( .A(n3003), .B(n2954), .Z(n3007) );
  OR2 U1305 ( .A(n3001), .B(n3002), .Z(n3006) );
  OR2 U1306 ( .A(n2999), .B(n3000), .Z(n3005) );
  OR2 U1307 ( .A(n2997), .B(n2998), .Z(n3004) );
  OR2 U1308 ( .A(n2995), .B(n2996), .Z(n3003) );
  OR2 U1309 ( .A(n2993), .B(n2994), .Z(n3002) );
  OR2 U1310 ( .A(n2991), .B(n2992), .Z(n3001) );
  OR2 U1311 ( .A(n2989), .B(n2990), .Z(n3000) );
  OR2 U1312 ( .A(n2987), .B(n2988), .Z(n2999) );
  OR2 U1313 ( .A(n2985), .B(n2986), .Z(n2998) );
  OR2 U1314 ( .A(n2983), .B(n2984), .Z(n2997) );
  OR2 U1315 ( .A(n2981), .B(n2982), .Z(n2996) );
  OR2 U1316 ( .A(n2979), .B(n2980), .Z(n2995) );
  OR2 U1317 ( .A(n2977), .B(n2978), .Z(n2994) );
  OR2 U1318 ( .A(n2975), .B(n2976), .Z(n2993) );
  OR2 U1319 ( .A(n2973), .B(n2974), .Z(n2992) );
  OR2 U1320 ( .A(n2971), .B(n2972), .Z(n2991) );
  OR2 U1321 ( .A(n2969), .B(n2970), .Z(n2990) );
  OR2 U1322 ( .A(n2967), .B(n2968), .Z(n2989) );
  OR2 U1323 ( .A(n2965), .B(n2966), .Z(n2988) );
  OR2 U1324 ( .A(n2963), .B(n2964), .Z(n2987) );
  OR2 U1325 ( .A(n2961), .B(n2962), .Z(n2986) );
  OR2 U1326 ( .A(n2959), .B(n2960), .Z(n2985) );
  OR2 U1327 ( .A(n2957), .B(n2958), .Z(n2984) );
  OR2 U1328 ( .A(n2955), .B(n2956), .Z(n2983) );
  OR2 U1329 ( .A(n2952), .B(n2953), .Z(n2982) );
  OR2 U1330 ( .A(n2950), .B(n2951), .Z(n2981) );
  OR2 U1331 ( .A(n2948), .B(n2949), .Z(n2980) );
  OR2 U1332 ( .A(n2946), .B(n2947), .Z(n2979) );
  OR2 U1333 ( .A(n2944), .B(n2945), .Z(n2978) );
  OR2 U1334 ( .A(n2942), .B(n2943), .Z(n2977) );
  OR2 U1335 ( .A(n2940), .B(n2941), .Z(n2976) );
  OR2 U1336 ( .A(n2938), .B(n2939), .Z(n2975) );
  OR2 U1337 ( .A(n2936), .B(n2937), .Z(n2974) );
  OR2 U1338 ( .A(n2934), .B(n2935), .Z(n2973) );
  OR2 U1339 ( .A(n2932), .B(n2933), .Z(n2972) );
  OR2 U1340 ( .A(n2930), .B(n2931), .Z(n2971) );
  OR2 U1341 ( .A(n2928), .B(n2929), .Z(n2970) );
  OR2 U1342 ( .A(n2926), .B(n2927), .Z(n2969) );
  OR2 U1343 ( .A(n2924), .B(n2925), .Z(n2968) );
  OR2 U1344 ( .A(n2922), .B(n2923), .Z(n2967) );
  OR2 U1345 ( .A(n2920), .B(n2921), .Z(n2966) );
  OR2 U1346 ( .A(n2918), .B(n2919), .Z(n2965) );
  OR2 U1347 ( .A(n2916), .B(n2917), .Z(n2964) );
  OR2 U1348 ( .A(n2914), .B(n2915), .Z(n2963) );
  OR2 U1349 ( .A(n2912), .B(n2913), .Z(n2962) );
  OR2 U1350 ( .A(n2910), .B(n2911), .Z(n2961) );
  OR2 U1351 ( .A(n2908), .B(n2909), .Z(n2960) );
  OR2 U1352 ( .A(n2906), .B(n2907), .Z(n2959) );
  OR2 U1353 ( .A(n2904), .B(n2905), .Z(n2958) );
  OR2 U1354 ( .A(n2902), .B(n2903), .Z(n2957) );
  OR2 U1355 ( .A(n2790), .B(n2901), .Z(n2956) );
  OR2 U1356 ( .A(n2899), .B(n2900), .Z(n2955) );
  OR2 U1357 ( .A(n2897), .B(n2898), .Z(n2954) );
  OR2 U1358 ( .A(n2895), .B(n2896), .Z(n2953) );
  OR2 U1359 ( .A(n2893), .B(n2894), .Z(n2952) );
  OR2 U1360 ( .A(n2891), .B(n2892), .Z(n2951) );
  OR2 U1361 ( .A(n2889), .B(n2890), .Z(n2950) );
  OR2 U1362 ( .A(n2887), .B(n2888), .Z(n2949) );
  OR2 U1363 ( .A(n2885), .B(n2886), .Z(n2948) );
  OR2 U1364 ( .A(n2883), .B(n2884), .Z(n2947) );
  OR2 U1365 ( .A(n2881), .B(n2882), .Z(n2946) );
  OR2 U1366 ( .A(n2879), .B(n2880), .Z(n2945) );
  OR2 U1367 ( .A(n2877), .B(n2878), .Z(n2944) );
  OR2 U1368 ( .A(n2875), .B(n2876), .Z(n2943) );
  OR2 U1369 ( .A(n2873), .B(n2874), .Z(n2942) );
  OR2 U1370 ( .A(n2871), .B(n2872), .Z(n2941) );
  OR2 U1371 ( .A(n2869), .B(n2870), .Z(n2940) );
  OR2 U1372 ( .A(n2867), .B(n2868), .Z(n2939) );
  OR2 U1373 ( .A(n2865), .B(n2866), .Z(n2938) );
  OR2 U1374 ( .A(n2863), .B(n2864), .Z(n2937) );
  OR2 U1375 ( .A(n2861), .B(n2862), .Z(n2936) );
  OR2 U1376 ( .A(n2859), .B(n2860), .Z(n2935) );
  OR2 U1377 ( .A(n2857), .B(n2858), .Z(n2934) );
  OR2 U1378 ( .A(n2855), .B(n2856), .Z(n2933) );
  OR2 U1379 ( .A(n2853), .B(n2854), .Z(n2932) );
  OR2 U1380 ( .A(n2851), .B(n2852), .Z(n2931) );
  OR2 U1381 ( .A(n2849), .B(n2850), .Z(n2930) );
  OR2 U1382 ( .A(n2847), .B(n2848), .Z(n2929) );
  OR2 U1383 ( .A(n2845), .B(n2846), .Z(n2928) );
  OR2 U1384 ( .A(n2843), .B(n2844), .Z(n2927) );
  OR2 U1385 ( .A(n2841), .B(n2842), .Z(n2926) );
  OR2 U1386 ( .A(n2839), .B(n2840), .Z(n2925) );
  OR2 U1387 ( .A(n2837), .B(n2838), .Z(n2924) );
  OR2 U1388 ( .A(n2835), .B(n2836), .Z(n2923) );
  OR2 U1389 ( .A(n2833), .B(n2834), .Z(n2922) );
  OR2 U1390 ( .A(n2831), .B(n2832), .Z(n2921) );
  OR2 U1391 ( .A(n2829), .B(n2830), .Z(n2920) );
  OR2 U1392 ( .A(n2827), .B(n2828), .Z(n2919) );
  OR2 U1393 ( .A(n2825), .B(n2826), .Z(n2918) );
  OR2 U1394 ( .A(n2823), .B(n2824), .Z(n2917) );
  OR2 U1395 ( .A(n2821), .B(n2822), .Z(n2916) );
  OR2 U1396 ( .A(n2819), .B(n2820), .Z(n2915) );
  OR2 U1397 ( .A(n2817), .B(n2818), .Z(n2914) );
  OR2 U1398 ( .A(n2815), .B(n2816), .Z(n2913) );
  OR2 U1399 ( .A(n2813), .B(n2814), .Z(n2912) );
  OR2 U1400 ( .A(n2811), .B(n2812), .Z(n2911) );
  OR2 U1401 ( .A(n2809), .B(n2810), .Z(n2910) );
  OR2 U1402 ( .A(n2807), .B(n2808), .Z(n2909) );
  OR2 U1403 ( .A(n2805), .B(n2806), .Z(n2908) );
  OR2 U1404 ( .A(n2803), .B(n2804), .Z(n2907) );
  OR2 U1405 ( .A(n2801), .B(n2802), .Z(n2906) );
  OR2 U1406 ( .A(n2799), .B(n2800), .Z(n2905) );
  OR2 U1407 ( .A(n2797), .B(n2798), .Z(n2904) );
  OR2 U1408 ( .A(n2795), .B(n2796), .Z(n2903) );
  OR2 U1409 ( .A(n2793), .B(n2794), .Z(n2902) );
  OR2 U1410 ( .A(n2791), .B(n2792), .Z(n2901) );
  OR2 U1411 ( .A(n2789), .B(N1120), .Z(n2900) );
  OR2 U1412 ( .A(n2787), .B(n2788), .Z(n2899) );
  AN2 U1413 ( .A(pos_disp_tx), .B(N8311), .Z(n2898) );
  AN2 U1414 ( .A(n291), .B(n153), .Z(n2897) );
  AN2 U1415 ( .A(pos_disp_tx), .B(n33), .Z(n2896) );
  AN2 U1416 ( .A(n291), .B(n19), .Z(n2895) );
  AN2 U1417 ( .A(n291), .B(n172), .Z(n2894) );
  AN2 U1418 ( .A(n291), .B(n26), .Z(n2893) );
  AN2 U1419 ( .A(n291), .B(n178), .Z(n2892) );
  AN2 U1420 ( .A(n291), .B(n23), .Z(n2891) );
  AN2 U1421 ( .A(n291), .B(n173), .Z(n2890) );
  AN2 U1422 ( .A(n291), .B(n27), .Z(n2889) );
  AN2 U1423 ( .A(n291), .B(n176), .Z(n2888) );
  AN2 U1424 ( .A(pos_disp_tx), .B(n166), .Z(n2887) );
  AN2 U1425 ( .A(n291), .B(n44), .Z(n2886) );
  AN2 U1426 ( .A(pos_disp_tx), .B(n179), .Z(n2885) );
  AN2 U1427 ( .A(pos_disp_tx), .B(n24), .Z(n2884) );
  AN2 U1428 ( .A(n291), .B(n155), .Z(n2883) );
  AN2 U1429 ( .A(pos_disp_tx), .B(n35), .Z(n2882) );
  AN2 U1430 ( .A(n291), .B(n21), .Z(n2881) );
  AN2 U1431 ( .A(n291), .B(n174), .Z(n2880) );
  AN2 U1432 ( .A(n291), .B(n28), .Z(n2879) );
  AN2 U1433 ( .A(n291), .B(n180), .Z(n2878) );
  AN2 U1434 ( .A(n291), .B(n25), .Z(n2877) );
  AN2 U1435 ( .A(n291), .B(n205), .Z(n2876) );
  AN2 U1436 ( .A(n291), .B(n29), .Z(n2875) );
  AN2 U1437 ( .A(n291), .B(n218), .Z(n2874) );
  AN2 U1438 ( .A(pos_disp_tx), .B(n267), .Z(n2873) );
  AN2 U1439 ( .A(n291), .B(n133), .Z(n2872) );
  AN2 U1440 ( .A(pos_disp_tx), .B(n181), .Z(n2871) );
  AN2 U1441 ( .A(pos_disp_tx), .B(n60), .Z(n2870) );
  AN2 U1442 ( .A(n291), .B(n231), .Z(n2869) );
  AN2 U1443 ( .A(pos_disp_tx), .B(n97), .Z(n2868) );
  AN2 U1444 ( .A(n291), .B(n48), .Z(n2867) );
  AN2 U1445 ( .A(n291), .B(n206), .Z(n2866) );
  AN2 U1446 ( .A(n291), .B(n72), .Z(n2865) );
  AN2 U1447 ( .A(n291), .B(n182), .Z(n2864) );
  AN2 U1448 ( .A(n291), .B(n61), .Z(n2863) );
  AN2 U1449 ( .A(n291), .B(n207), .Z(n2862) );
  AN2 U1450 ( .A(n291), .B(n73), .Z(n2861) );
  AN2 U1451 ( .A(n291), .B(n220), .Z(n2860) );
  AN2 U1452 ( .A(pos_disp_tx), .B(n269), .Z(n2859) );
  AN2 U1453 ( .A(n291), .B(n135), .Z(n2858) );
  AN2 U1454 ( .A(pos_disp_tx), .B(n183), .Z(n2857) );
  AN2 U1455 ( .A(pos_disp_tx), .B(n62), .Z(n2856) );
  AN2 U1456 ( .A(n291), .B(n233), .Z(n2855) );
  AN2 U1457 ( .A(pos_disp_tx), .B(n99), .Z(n2854) );
  AN2 U1458 ( .A(n291), .B(n50), .Z(n2853) );
  AN2 U1459 ( .A(n291), .B(n208), .Z(n2852) );
  AN2 U1460 ( .A(n291), .B(n74), .Z(n2851) );
  AN2 U1461 ( .A(n291), .B(n184), .Z(n2850) );
  AN2 U1462 ( .A(n291), .B(n63), .Z(n2849) );
  AN2 U1463 ( .A(n291), .B(n209), .Z(n2848) );
  AN2 U1464 ( .A(n291), .B(n75), .Z(n2847) );
  AN2 U1465 ( .A(n291), .B(n222), .Z(n2846) );
  AN2 U1466 ( .A(pos_disp_tx), .B(n271), .Z(n2845) );
  AN2 U1467 ( .A(n291), .B(n137), .Z(n2844) );
  AN2 U1468 ( .A(pos_disp_tx), .B(n185), .Z(n2843) );
  AN2 U1469 ( .A(pos_disp_tx), .B(n64), .Z(n2842) );
  AN2 U1470 ( .A(n291), .B(n235), .Z(n2841) );
  AN2 U1471 ( .A(pos_disp_tx), .B(n101), .Z(n2840) );
  AN2 U1472 ( .A(n291), .B(n52), .Z(n2839) );
  AN2 U1473 ( .A(n291), .B(n210), .Z(n2838) );
  AN2 U1474 ( .A(n291), .B(n76), .Z(n2837) );
  AN2 U1475 ( .A(n291), .B(n186), .Z(n2836) );
  AN2 U1476 ( .A(n291), .B(n65), .Z(n2835) );
  AN2 U1477 ( .A(n291), .B(n211), .Z(n2834) );
  AN2 U1478 ( .A(n291), .B(n77), .Z(n2833) );
  AN2 U1479 ( .A(n291), .B(n224), .Z(n2832) );
  AN2 U1480 ( .A(pos_disp_tx), .B(n273), .Z(n2831) );
  AN2 U1481 ( .A(n291), .B(n139), .Z(n2830) );
  AN2 U1482 ( .A(pos_disp_tx), .B(n187), .Z(n2829) );
  AN2 U1483 ( .A(pos_disp_tx), .B(n66), .Z(n2828) );
  AN2 U1484 ( .A(n291), .B(n237), .Z(n2827) );
  AN2 U1485 ( .A(pos_disp_tx), .B(n103), .Z(n2826) );
  AN2 U1486 ( .A(n291), .B(n54), .Z(n2825) );
  AN2 U1487 ( .A(n291), .B(n212), .Z(n2824) );
  AN2 U1488 ( .A(n291), .B(n78), .Z(n2823) );
  AN2 U1489 ( .A(n291), .B(n188), .Z(n2822) );
  AN2 U1490 ( .A(n291), .B(n67), .Z(n2821) );
  AN2 U1491 ( .A(n291), .B(n213), .Z(n2820) );
  AN2 U1492 ( .A(n291), .B(n79), .Z(n2819) );
  AN2 U1493 ( .A(n291), .B(n226), .Z(n2818) );
  AN2 U1494 ( .A(pos_disp_tx), .B(n275), .Z(n2817) );
  AN2 U1495 ( .A(n291), .B(n141), .Z(n2816) );
  AN2 U1496 ( .A(pos_disp_tx), .B(n189), .Z(n2815) );
  AN2 U1497 ( .A(pos_disp_tx), .B(n68), .Z(n2814) );
  AN2 U1498 ( .A(n291), .B(n239), .Z(n2813) );
  AN2 U1499 ( .A(pos_disp_tx), .B(n105), .Z(n2812) );
  AN2 U1500 ( .A(n291), .B(n56), .Z(n2811) );
  AN2 U1501 ( .A(n291), .B(n214), .Z(n2810) );
  AN2 U1502 ( .A(n291), .B(n80), .Z(n2809) );
  AN2 U1503 ( .A(n291), .B(n190), .Z(n2808) );
  AN2 U1504 ( .A(n291), .B(n69), .Z(n2807) );
  AN2 U1505 ( .A(n291), .B(n215), .Z(n2806) );
  AN2 U1506 ( .A(n291), .B(n81), .Z(n2805) );
  AN2 U1507 ( .A(n291), .B(n228), .Z(n2804) );
  AN2 U1508 ( .A(pos_disp_tx), .B(n277), .Z(n2803) );
  AN2 U1509 ( .A(n291), .B(n143), .Z(n2802) );
  AN2 U1510 ( .A(pos_disp_tx), .B(n191), .Z(n2801) );
  AN2 U1511 ( .A(pos_disp_tx), .B(n70), .Z(n2800) );
  AN2 U1512 ( .A(n291), .B(n241), .Z(n2799) );
  AN2 U1513 ( .A(pos_disp_tx), .B(n107), .Z(n2798) );
  AN2 U1514 ( .A(n291), .B(n58), .Z(n2797) );
  AN2 U1515 ( .A(n291), .B(n216), .Z(n2796) );
  AN2 U1516 ( .A(n291), .B(n82), .Z(n2795) );
  AN2 U1517 ( .A(n291), .B(n192), .Z(n2794) );
  AN2 U1518 ( .A(n291), .B(n71), .Z(n2793) );
  AN2 U1519 ( .A(n291), .B(n217), .Z(n2792) );
  AN2 U1520 ( .A(n291), .B(n83), .Z(n2791) );
  AN2 U1521 ( .A(n291), .B(n230), .Z(n2790) );
  AN2 U1522 ( .A(pos_disp_tx), .B(n279), .Z(n2789) );
  AN2 U1523 ( .A(n291), .B(n145), .Z(n2788) );
  AN2 U1524 ( .A(pos_disp_tx), .B(N239), .Z(n2787) );
  OR2 U1525 ( .A(n2785), .B(n2786), .Z(N839) );
  OR2 U1526 ( .A(n2783), .B(n2784), .Z(n2786) );
  OR2 U1527 ( .A(n2781), .B(n2782), .Z(n2785) );
  OR2 U1528 ( .A(n2780), .B(n2731), .Z(n2784) );
  OR2 U1529 ( .A(n2778), .B(n2779), .Z(n2783) );
  OR2 U1530 ( .A(n2776), .B(n2777), .Z(n2782) );
  OR2 U1531 ( .A(n2774), .B(n2775), .Z(n2781) );
  OR2 U1532 ( .A(n2772), .B(n2773), .Z(n2780) );
  OR2 U1533 ( .A(n2770), .B(n2771), .Z(n2779) );
  OR2 U1534 ( .A(n2768), .B(n2769), .Z(n2778) );
  OR2 U1535 ( .A(n2766), .B(n2767), .Z(n2777) );
  OR2 U1536 ( .A(n2764), .B(n2765), .Z(n2776) );
  OR2 U1537 ( .A(n2762), .B(n2763), .Z(n2775) );
  OR2 U1538 ( .A(n2760), .B(n2761), .Z(n2774) );
  OR2 U1539 ( .A(n2758), .B(n2759), .Z(n2773) );
  OR2 U1540 ( .A(n2756), .B(n2757), .Z(n2772) );
  OR2 U1541 ( .A(n2754), .B(n2755), .Z(n2771) );
  OR2 U1542 ( .A(n2752), .B(n2753), .Z(n2770) );
  OR2 U1543 ( .A(n2750), .B(n2751), .Z(n2769) );
  OR2 U1544 ( .A(n2748), .B(n2749), .Z(n2768) );
  OR2 U1545 ( .A(n2746), .B(n2747), .Z(n2767) );
  OR2 U1546 ( .A(n2744), .B(n2745), .Z(n2766) );
  OR2 U1547 ( .A(n2742), .B(n2743), .Z(n2765) );
  OR2 U1548 ( .A(n2740), .B(n2741), .Z(n2764) );
  OR2 U1549 ( .A(n2738), .B(n2739), .Z(n2763) );
  OR2 U1550 ( .A(n2736), .B(n2737), .Z(n2762) );
  OR2 U1551 ( .A(n2734), .B(n2735), .Z(n2761) );
  OR2 U1552 ( .A(n2732), .B(n2733), .Z(n2760) );
  OR2 U1553 ( .A(n2729), .B(n2730), .Z(n2759) );
  OR2 U1554 ( .A(n2727), .B(n2728), .Z(n2758) );
  OR2 U1555 ( .A(n2725), .B(n2726), .Z(n2757) );
  OR2 U1556 ( .A(n2723), .B(n2724), .Z(n2756) );
  OR2 U1557 ( .A(n2721), .B(n2722), .Z(n2755) );
  OR2 U1558 ( .A(n2719), .B(n2720), .Z(n2754) );
  OR2 U1559 ( .A(n2717), .B(n2718), .Z(n2753) );
  OR2 U1560 ( .A(n2715), .B(n2716), .Z(n2752) );
  OR2 U1561 ( .A(n2713), .B(n2714), .Z(n2751) );
  OR2 U1562 ( .A(n2711), .B(n2712), .Z(n2750) );
  OR2 U1563 ( .A(n2709), .B(n2710), .Z(n2749) );
  OR2 U1564 ( .A(n2707), .B(n2708), .Z(n2748) );
  OR2 U1565 ( .A(n2705), .B(n2706), .Z(n2747) );
  OR2 U1566 ( .A(n2703), .B(n2704), .Z(n2746) );
  OR2 U1567 ( .A(n2701), .B(n2702), .Z(n2745) );
  OR2 U1568 ( .A(n2699), .B(n2700), .Z(n2744) );
  OR2 U1569 ( .A(n2697), .B(n2698), .Z(n2743) );
  OR2 U1570 ( .A(n2695), .B(n2696), .Z(n2742) );
  OR2 U1571 ( .A(n2693), .B(n2694), .Z(n2741) );
  OR2 U1572 ( .A(n2691), .B(n2692), .Z(n2740) );
  OR2 U1573 ( .A(n2689), .B(n2690), .Z(n2739) );
  OR2 U1574 ( .A(n2687), .B(n2688), .Z(n2738) );
  OR2 U1575 ( .A(n2685), .B(n2686), .Z(n2737) );
  OR2 U1576 ( .A(n2683), .B(n2684), .Z(n2736) );
  OR2 U1577 ( .A(n2681), .B(n2682), .Z(n2735) );
  OR2 U1578 ( .A(n2679), .B(n2680), .Z(n2734) );
  OR2 U1579 ( .A(n2677), .B(n2678), .Z(n2733) );
  OR2 U1580 ( .A(n2676), .B(n2566), .Z(n2732) );
  OR2 U1581 ( .A(n2674), .B(n2675), .Z(n2731) );
  OR2 U1582 ( .A(n2672), .B(n2673), .Z(n2730) );
  OR2 U1583 ( .A(n2670), .B(n2671), .Z(n2729) );
  OR2 U1584 ( .A(n2668), .B(n2669), .Z(n2728) );
  OR2 U1585 ( .A(n2666), .B(n2667), .Z(n2727) );
  OR2 U1586 ( .A(n2664), .B(n2665), .Z(n2726) );
  OR2 U1587 ( .A(n2662), .B(n2663), .Z(n2725) );
  OR2 U1588 ( .A(n2660), .B(n2661), .Z(n2724) );
  OR2 U1589 ( .A(n2658), .B(n2659), .Z(n2723) );
  OR2 U1590 ( .A(n2656), .B(n2657), .Z(n2722) );
  OR2 U1591 ( .A(n2654), .B(n2655), .Z(n2721) );
  OR2 U1592 ( .A(n2652), .B(n2653), .Z(n2720) );
  OR2 U1593 ( .A(n2650), .B(n2651), .Z(n2719) );
  OR2 U1594 ( .A(n2648), .B(n2649), .Z(n2718) );
  OR2 U1595 ( .A(n2646), .B(n2647), .Z(n2717) );
  OR2 U1596 ( .A(n2644), .B(n2645), .Z(n2716) );
  OR2 U1597 ( .A(n2642), .B(n2643), .Z(n2715) );
  OR2 U1598 ( .A(n2640), .B(n2641), .Z(n2714) );
  OR2 U1599 ( .A(n2638), .B(n2639), .Z(n2713) );
  OR2 U1600 ( .A(n2636), .B(n2637), .Z(n2712) );
  OR2 U1601 ( .A(n2634), .B(n2635), .Z(n2711) );
  OR2 U1602 ( .A(n2632), .B(n2633), .Z(n2710) );
  OR2 U1603 ( .A(n2630), .B(n2631), .Z(n2709) );
  OR2 U1604 ( .A(n2628), .B(n2629), .Z(n2708) );
  OR2 U1605 ( .A(n2626), .B(n2627), .Z(n2707) );
  OR2 U1606 ( .A(n2624), .B(n2625), .Z(n2706) );
  OR2 U1607 ( .A(n2622), .B(n2623), .Z(n2705) );
  OR2 U1608 ( .A(n2620), .B(n2621), .Z(n2704) );
  OR2 U1609 ( .A(n2618), .B(n2619), .Z(n2703) );
  OR2 U1610 ( .A(n2616), .B(n2617), .Z(n2702) );
  OR2 U1611 ( .A(n2614), .B(n2615), .Z(n2701) );
  OR2 U1612 ( .A(n2612), .B(n2613), .Z(n2700) );
  OR2 U1613 ( .A(n2610), .B(n2611), .Z(n2699) );
  OR2 U1614 ( .A(n2608), .B(n2609), .Z(n2698) );
  OR2 U1615 ( .A(n2606), .B(n2607), .Z(n2697) );
  OR2 U1616 ( .A(n2604), .B(n2605), .Z(n2696) );
  OR2 U1617 ( .A(n2602), .B(n2603), .Z(n2695) );
  OR2 U1618 ( .A(n2600), .B(n2601), .Z(n2694) );
  OR2 U1619 ( .A(n2598), .B(n2599), .Z(n2693) );
  OR2 U1620 ( .A(n2596), .B(n2597), .Z(n2692) );
  OR2 U1621 ( .A(n2594), .B(n2595), .Z(n2691) );
  OR2 U1622 ( .A(n2592), .B(n2593), .Z(n2690) );
  OR2 U1623 ( .A(n2590), .B(n2591), .Z(n2689) );
  OR2 U1624 ( .A(n2588), .B(n2589), .Z(n2688) );
  OR2 U1625 ( .A(n2586), .B(n2587), .Z(n2687) );
  OR2 U1626 ( .A(n2584), .B(n2585), .Z(n2686) );
  OR2 U1627 ( .A(n2582), .B(n2583), .Z(n2685) );
  OR2 U1628 ( .A(n2580), .B(n2581), .Z(n2684) );
  OR2 U1629 ( .A(n2578), .B(n2579), .Z(n2683) );
  OR2 U1630 ( .A(n2576), .B(n2577), .Z(n2682) );
  OR2 U1631 ( .A(n2574), .B(n2575), .Z(n2681) );
  OR2 U1632 ( .A(n2572), .B(n2573), .Z(n2680) );
  OR2 U1633 ( .A(n2570), .B(n2571), .Z(n2679) );
  OR2 U1634 ( .A(n2568), .B(n2569), .Z(n2678) );
  OR2 U1635 ( .A(n2567), .B(N11011), .Z(n2677) );
  OR2 U1636 ( .A(n2564), .B(n2565), .Z(n2676) );
  AN2 U1637 ( .A(n291), .B(N8311), .Z(n2675) );
  AN2 U1638 ( .A(n291), .B(n153), .Z(n2674) );
  AN2 U1639 ( .A(n291), .B(n33), .Z(n2673) );
  AN2 U1640 ( .A(pos_disp_tx), .B(n19), .Z(n2672) );
  AN2 U1641 ( .A(pos_disp_tx), .B(n172), .Z(n2671) );
  AN2 U1642 ( .A(n291), .B(n26), .Z(n2670) );
  AN2 U1643 ( .A(n291), .B(n178), .Z(n2669) );
  AN2 U1644 ( .A(pos_disp_tx), .B(n23), .Z(n2668) );
  AN2 U1645 ( .A(n291), .B(n173), .Z(n2667) );
  AN2 U1646 ( .A(n291), .B(n27), .Z(n2666) );
  AN2 U1647 ( .A(pos_disp_tx), .B(n176), .Z(n2665) );
  AN2 U1648 ( .A(n291), .B(n166), .Z(n2664) );
  AN2 U1649 ( .A(n291), .B(n44), .Z(n2663) );
  AN2 U1650 ( .A(pos_disp_tx), .B(n179), .Z(n2662) );
  AN2 U1651 ( .A(n291), .B(n24), .Z(n2661) );
  AN2 U1652 ( .A(n291), .B(n155), .Z(n2660) );
  AN2 U1653 ( .A(n291), .B(n35), .Z(n2659) );
  AN2 U1654 ( .A(pos_disp_tx), .B(n21), .Z(n2658) );
  AN2 U1655 ( .A(pos_disp_tx), .B(n174), .Z(n2657) );
  AN2 U1656 ( .A(n291), .B(n28), .Z(n2656) );
  AN2 U1657 ( .A(n291), .B(n180), .Z(n2655) );
  AN2 U1658 ( .A(pos_disp_tx), .B(n25), .Z(n2654) );
  AN2 U1659 ( .A(n291), .B(n205), .Z(n2653) );
  AN2 U1660 ( .A(n291), .B(n29), .Z(n2652) );
  AN2 U1661 ( .A(pos_disp_tx), .B(n218), .Z(n2651) );
  AN2 U1662 ( .A(n291), .B(n267), .Z(n2650) );
  AN2 U1663 ( .A(n291), .B(n133), .Z(n2649) );
  AN2 U1664 ( .A(pos_disp_tx), .B(n181), .Z(n2648) );
  AN2 U1665 ( .A(n291), .B(n60), .Z(n2647) );
  AN2 U1666 ( .A(n291), .B(n231), .Z(n2646) );
  AN2 U1667 ( .A(n291), .B(n97), .Z(n2645) );
  AN2 U1668 ( .A(pos_disp_tx), .B(n48), .Z(n2644) );
  AN2 U1669 ( .A(pos_disp_tx), .B(n206), .Z(n2643) );
  AN2 U1670 ( .A(n291), .B(n72), .Z(n2642) );
  AN2 U1671 ( .A(n291), .B(n182), .Z(n2641) );
  AN2 U1672 ( .A(pos_disp_tx), .B(n61), .Z(n2640) );
  AN2 U1673 ( .A(n291), .B(n207), .Z(n2639) );
  AN2 U1674 ( .A(n291), .B(n73), .Z(n2638) );
  AN2 U1675 ( .A(pos_disp_tx), .B(n220), .Z(n2637) );
  AN2 U1676 ( .A(n291), .B(n269), .Z(n2636) );
  AN2 U1677 ( .A(n291), .B(n135), .Z(n2635) );
  AN2 U1678 ( .A(pos_disp_tx), .B(n183), .Z(n2634) );
  AN2 U1679 ( .A(n291), .B(n62), .Z(n2633) );
  AN2 U1680 ( .A(n291), .B(n233), .Z(n2632) );
  AN2 U1681 ( .A(n291), .B(n99), .Z(n2631) );
  AN2 U1682 ( .A(pos_disp_tx), .B(n50), .Z(n2630) );
  AN2 U1683 ( .A(pos_disp_tx), .B(n208), .Z(n2629) );
  AN2 U1684 ( .A(n291), .B(n74), .Z(n2628) );
  AN2 U1685 ( .A(n291), .B(n184), .Z(n2627) );
  AN2 U1686 ( .A(pos_disp_tx), .B(n63), .Z(n2626) );
  AN2 U1687 ( .A(n291), .B(n209), .Z(n2625) );
  AN2 U1688 ( .A(n291), .B(n75), .Z(n2624) );
  AN2 U1689 ( .A(pos_disp_tx), .B(n222), .Z(n2623) );
  AN2 U1690 ( .A(n291), .B(n271), .Z(n2622) );
  AN2 U1691 ( .A(n291), .B(n137), .Z(n2621) );
  AN2 U1692 ( .A(pos_disp_tx), .B(n185), .Z(n2620) );
  AN2 U1693 ( .A(n291), .B(n64), .Z(n2619) );
  AN2 U1694 ( .A(n291), .B(n235), .Z(n2618) );
  AN2 U1695 ( .A(n291), .B(n101), .Z(n2617) );
  AN2 U1696 ( .A(pos_disp_tx), .B(n52), .Z(n2616) );
  AN2 U1697 ( .A(pos_disp_tx), .B(n210), .Z(n2615) );
  AN2 U1698 ( .A(n291), .B(n76), .Z(n2614) );
  AN2 U1699 ( .A(n291), .B(n186), .Z(n2613) );
  AN2 U1700 ( .A(pos_disp_tx), .B(n65), .Z(n2612) );
  AN2 U1701 ( .A(n291), .B(n211), .Z(n2611) );
  AN2 U1702 ( .A(n291), .B(n77), .Z(n2610) );
  AN2 U1703 ( .A(pos_disp_tx), .B(n224), .Z(n2609) );
  AN2 U1704 ( .A(n291), .B(n273), .Z(n2608) );
  AN2 U1705 ( .A(n291), .B(n139), .Z(n2607) );
  AN2 U1706 ( .A(pos_disp_tx), .B(n187), .Z(n2606) );
  AN2 U1707 ( .A(n291), .B(n66), .Z(n2605) );
  AN2 U1708 ( .A(n291), .B(n237), .Z(n2604) );
  AN2 U1709 ( .A(n291), .B(n103), .Z(n2603) );
  AN2 U1710 ( .A(pos_disp_tx), .B(n54), .Z(n2602) );
  AN2 U1711 ( .A(pos_disp_tx), .B(n212), .Z(n2601) );
  AN2 U1712 ( .A(n291), .B(n78), .Z(n2600) );
  AN2 U1713 ( .A(n291), .B(n188), .Z(n2599) );
  AN2 U1714 ( .A(pos_disp_tx), .B(n67), .Z(n2598) );
  AN2 U1715 ( .A(n291), .B(n213), .Z(n2597) );
  AN2 U1716 ( .A(n291), .B(n79), .Z(n2596) );
  AN2 U1717 ( .A(pos_disp_tx), .B(n226), .Z(n2595) );
  AN2 U1718 ( .A(n291), .B(n275), .Z(n2594) );
  AN2 U1719 ( .A(n291), .B(n141), .Z(n2593) );
  AN2 U1720 ( .A(pos_disp_tx), .B(n189), .Z(n2592) );
  AN2 U1721 ( .A(n291), .B(n68), .Z(n2591) );
  AN2 U1722 ( .A(n291), .B(n239), .Z(n2590) );
  AN2 U1723 ( .A(n291), .B(n105), .Z(n2589) );
  AN2 U1724 ( .A(pos_disp_tx), .B(n56), .Z(n2588) );
  AN2 U1725 ( .A(pos_disp_tx), .B(n214), .Z(n2587) );
  AN2 U1726 ( .A(n291), .B(n80), .Z(n2586) );
  AN2 U1727 ( .A(n291), .B(n190), .Z(n2585) );
  AN2 U1728 ( .A(pos_disp_tx), .B(n69), .Z(n2584) );
  AN2 U1729 ( .A(n291), .B(n215), .Z(n2583) );
  AN2 U1730 ( .A(n291), .B(n81), .Z(n2582) );
  AN2 U1731 ( .A(pos_disp_tx), .B(n228), .Z(n2581) );
  AN2 U1732 ( .A(n291), .B(n277), .Z(n2580) );
  AN2 U1733 ( .A(n291), .B(n143), .Z(n2579) );
  AN2 U1734 ( .A(pos_disp_tx), .B(n191), .Z(n2578) );
  AN2 U1735 ( .A(n291), .B(n70), .Z(n2577) );
  AN2 U1736 ( .A(n291), .B(n241), .Z(n2576) );
  AN2 U1737 ( .A(n291), .B(n107), .Z(n2575) );
  AN2 U1738 ( .A(pos_disp_tx), .B(n58), .Z(n2574) );
  AN2 U1739 ( .A(pos_disp_tx), .B(n216), .Z(n2573) );
  AN2 U1740 ( .A(n291), .B(n82), .Z(n2572) );
  AN2 U1741 ( .A(n291), .B(n192), .Z(n2571) );
  AN2 U1742 ( .A(pos_disp_tx), .B(n71), .Z(n2570) );
  AN2 U1743 ( .A(n291), .B(n217), .Z(n2569) );
  AN2 U1744 ( .A(n291), .B(n83), .Z(n2568) );
  AN2 U1745 ( .A(pos_disp_tx), .B(n230), .Z(n2567) );
  AN2 U1746 ( .A(n291), .B(n279), .Z(n2566) );
  AN2 U1747 ( .A(n291), .B(n145), .Z(n2565) );
  AN2 U1748 ( .A(pos_disp_tx), .B(N239), .Z(n2564) );
  OR2 U1749 ( .A(n2562), .B(n2563), .Z(N838) );
  OR2 U1750 ( .A(n2560), .B(n2561), .Z(n2563) );
  OR2 U1751 ( .A(n2558), .B(n2559), .Z(n2562) );
  OR2 U1752 ( .A(n2557), .B(n2508), .Z(n2561) );
  OR2 U1753 ( .A(n2555), .B(n2556), .Z(n2560) );
  OR2 U1754 ( .A(n2553), .B(n2554), .Z(n2559) );
  OR2 U1755 ( .A(n2551), .B(n2552), .Z(n2558) );
  OR2 U1756 ( .A(n2549), .B(n2550), .Z(n2557) );
  OR2 U1757 ( .A(n2547), .B(n2548), .Z(n2556) );
  OR2 U1758 ( .A(n2545), .B(n2546), .Z(n2555) );
  OR2 U1759 ( .A(n2543), .B(n2544), .Z(n2554) );
  OR2 U1760 ( .A(n2541), .B(n2542), .Z(n2553) );
  OR2 U1761 ( .A(n2539), .B(n2540), .Z(n2552) );
  OR2 U1762 ( .A(n2537), .B(n2538), .Z(n2551) );
  OR2 U1763 ( .A(n2535), .B(n2536), .Z(n2550) );
  OR2 U1764 ( .A(n2533), .B(n2534), .Z(n2549) );
  OR2 U1765 ( .A(n2531), .B(n2532), .Z(n2548) );
  OR2 U1766 ( .A(n2529), .B(n2530), .Z(n2547) );
  OR2 U1767 ( .A(n2527), .B(n2528), .Z(n2546) );
  OR2 U1768 ( .A(n2525), .B(n2526), .Z(n2545) );
  OR2 U1769 ( .A(n2523), .B(n2524), .Z(n2544) );
  OR2 U1770 ( .A(n2521), .B(n2522), .Z(n2543) );
  OR2 U1771 ( .A(n2519), .B(n2520), .Z(n2542) );
  OR2 U1772 ( .A(n2517), .B(n2518), .Z(n2541) );
  OR2 U1773 ( .A(n2515), .B(n2516), .Z(n2540) );
  OR2 U1774 ( .A(n2513), .B(n2514), .Z(n2539) );
  OR2 U1775 ( .A(n2511), .B(n2512), .Z(n2538) );
  OR2 U1776 ( .A(n2509), .B(n2510), .Z(n2537) );
  OR2 U1777 ( .A(n2506), .B(n2507), .Z(n2536) );
  OR2 U1778 ( .A(n2504), .B(n2505), .Z(n2535) );
  OR2 U1779 ( .A(n2502), .B(n2503), .Z(n2534) );
  OR2 U1780 ( .A(n2500), .B(n2501), .Z(n2533) );
  OR2 U1781 ( .A(n2498), .B(n2499), .Z(n2532) );
  OR2 U1782 ( .A(n2496), .B(n2497), .Z(n2531) );
  OR2 U1783 ( .A(n2494), .B(n2495), .Z(n2530) );
  OR2 U1784 ( .A(n2492), .B(n2493), .Z(n2529) );
  OR2 U1785 ( .A(n2490), .B(n2491), .Z(n2528) );
  OR2 U1786 ( .A(n2488), .B(n2489), .Z(n2527) );
  OR2 U1787 ( .A(n2486), .B(n2487), .Z(n2526) );
  OR2 U1788 ( .A(n2484), .B(n2485), .Z(n2525) );
  OR2 U1789 ( .A(n2482), .B(n2483), .Z(n2524) );
  OR2 U1790 ( .A(n2480), .B(n2481), .Z(n2523) );
  OR2 U1791 ( .A(n2478), .B(n2479), .Z(n2522) );
  OR2 U1792 ( .A(n2476), .B(n2477), .Z(n2521) );
  OR2 U1793 ( .A(n2474), .B(n2475), .Z(n2520) );
  OR2 U1794 ( .A(n2472), .B(n2473), .Z(n2519) );
  OR2 U1795 ( .A(n2470), .B(n2471), .Z(n2518) );
  OR2 U1796 ( .A(n2468), .B(n2469), .Z(n2517) );
  OR2 U1797 ( .A(n2466), .B(n2467), .Z(n2516) );
  OR2 U1798 ( .A(n2464), .B(n2465), .Z(n2515) );
  OR2 U1799 ( .A(n2462), .B(n2463), .Z(n2514) );
  OR2 U1800 ( .A(n2460), .B(n2461), .Z(n2513) );
  OR2 U1801 ( .A(n2458), .B(n2459), .Z(n2512) );
  OR2 U1802 ( .A(n2456), .B(n2457), .Z(n2511) );
  OR2 U1803 ( .A(n2454), .B(n2455), .Z(n2510) );
  OR2 U1804 ( .A(n2453), .B(n2343), .Z(n2509) );
  OR2 U1805 ( .A(n2451), .B(n2452), .Z(n2508) );
  OR2 U1806 ( .A(n2449), .B(n2450), .Z(n2507) );
  OR2 U1807 ( .A(n2447), .B(n2448), .Z(n2506) );
  OR2 U1808 ( .A(n2445), .B(n2446), .Z(n2505) );
  OR2 U1809 ( .A(n2443), .B(n2444), .Z(n2504) );
  OR2 U1810 ( .A(n2441), .B(n2442), .Z(n2503) );
  OR2 U1811 ( .A(n2439), .B(n2440), .Z(n2502) );
  OR2 U1812 ( .A(n2437), .B(n2438), .Z(n2501) );
  OR2 U1813 ( .A(n2435), .B(n2436), .Z(n2500) );
  OR2 U1814 ( .A(n2433), .B(n2434), .Z(n2499) );
  OR2 U1815 ( .A(n2431), .B(n2432), .Z(n2498) );
  OR2 U1816 ( .A(n2429), .B(n2430), .Z(n2497) );
  OR2 U1817 ( .A(n2427), .B(n2428), .Z(n2496) );
  OR2 U1818 ( .A(n2425), .B(n2426), .Z(n2495) );
  OR2 U1819 ( .A(n2423), .B(n2424), .Z(n2494) );
  OR2 U1820 ( .A(n2421), .B(n2422), .Z(n2493) );
  OR2 U1821 ( .A(n2419), .B(n2420), .Z(n2492) );
  OR2 U1822 ( .A(n2417), .B(n2418), .Z(n2491) );
  OR2 U1823 ( .A(n2415), .B(n2416), .Z(n2490) );
  OR2 U1824 ( .A(n2413), .B(n2414), .Z(n2489) );
  OR2 U1825 ( .A(n2411), .B(n2412), .Z(n2488) );
  OR2 U1826 ( .A(n2409), .B(n2410), .Z(n2487) );
  OR2 U1827 ( .A(n2407), .B(n2408), .Z(n2486) );
  OR2 U1828 ( .A(n2405), .B(n2406), .Z(n2485) );
  OR2 U1829 ( .A(n2403), .B(n2404), .Z(n2484) );
  OR2 U1830 ( .A(n2401), .B(n2402), .Z(n2483) );
  OR2 U1831 ( .A(n2399), .B(n2400), .Z(n2482) );
  OR2 U1832 ( .A(n2397), .B(n2398), .Z(n2481) );
  OR2 U1833 ( .A(n2395), .B(n2396), .Z(n2480) );
  OR2 U1834 ( .A(n2393), .B(n2394), .Z(n2479) );
  OR2 U1835 ( .A(n2391), .B(n2392), .Z(n2478) );
  OR2 U1836 ( .A(n2389), .B(n2390), .Z(n2477) );
  OR2 U1837 ( .A(n2387), .B(n2388), .Z(n2476) );
  OR2 U1838 ( .A(n2385), .B(n2386), .Z(n2475) );
  OR2 U1839 ( .A(n2383), .B(n2384), .Z(n2474) );
  OR2 U1840 ( .A(n2381), .B(n2382), .Z(n2473) );
  OR2 U1841 ( .A(n2379), .B(n2380), .Z(n2472) );
  OR2 U1842 ( .A(n2377), .B(n2378), .Z(n2471) );
  OR2 U1843 ( .A(n2375), .B(n2376), .Z(n2470) );
  OR2 U1844 ( .A(n2373), .B(n2374), .Z(n2469) );
  OR2 U1845 ( .A(n2371), .B(n2372), .Z(n2468) );
  OR2 U1846 ( .A(n2369), .B(n2370), .Z(n2467) );
  OR2 U1847 ( .A(n2367), .B(n2368), .Z(n2466) );
  OR2 U1848 ( .A(n2365), .B(n2366), .Z(n2465) );
  OR2 U1849 ( .A(n2363), .B(n2364), .Z(n2464) );
  OR2 U1850 ( .A(n2361), .B(n2362), .Z(n2463) );
  OR2 U1851 ( .A(n2359), .B(n2360), .Z(n2462) );
  OR2 U1852 ( .A(n2357), .B(n2358), .Z(n2461) );
  OR2 U1853 ( .A(n2355), .B(n2356), .Z(n2460) );
  OR2 U1854 ( .A(n2353), .B(n2354), .Z(n2459) );
  OR2 U1855 ( .A(n2351), .B(n2352), .Z(n2458) );
  OR2 U1856 ( .A(n2349), .B(n2350), .Z(n2457) );
  OR2 U1857 ( .A(n2347), .B(n2348), .Z(n2456) );
  OR2 U1858 ( .A(n2346), .B(N1063), .Z(n2455) );
  OR2 U1859 ( .A(n2344), .B(n2345), .Z(n2454) );
  OR2 U1860 ( .A(n2341), .B(n2342), .Z(n2453) );
  AN2 U1861 ( .A(pos_disp_tx), .B(N8311), .Z(n2452) );
  AN2 U1862 ( .A(n291), .B(n153), .Z(n2451) );
  AN2 U1863 ( .A(n291), .B(n33), .Z(n2450) );
  AN2 U1864 ( .A(n291), .B(n19), .Z(n2449) );
  AN2 U1865 ( .A(pos_disp_tx), .B(n172), .Z(n2448) );
  AN2 U1866 ( .A(pos_disp_tx), .B(n26), .Z(n2447) );
  AN2 U1867 ( .A(pos_disp_tx), .B(n178), .Z(n2446) );
  AN2 U1868 ( .A(n291), .B(n23), .Z(n2445) );
  AN2 U1869 ( .A(pos_disp_tx), .B(n173), .Z(n2444) );
  AN2 U1870 ( .A(pos_disp_tx), .B(n27), .Z(n2443) );
  AN2 U1871 ( .A(n291), .B(n176), .Z(n2442) );
  AN2 U1872 ( .A(n291), .B(n166), .Z(n2441) );
  AN2 U1873 ( .A(n291), .B(n44), .Z(n2440) );
  AN2 U1874 ( .A(n291), .B(n179), .Z(n2439) );
  AN2 U1875 ( .A(pos_disp_tx), .B(n24), .Z(n2438) );
  AN2 U1876 ( .A(n291), .B(n155), .Z(n2437) );
  AN2 U1877 ( .A(n291), .B(n35), .Z(n2436) );
  AN2 U1878 ( .A(n291), .B(n21), .Z(n2435) );
  AN2 U1879 ( .A(pos_disp_tx), .B(n174), .Z(n2434) );
  AN2 U1880 ( .A(pos_disp_tx), .B(n28), .Z(n2433) );
  AN2 U1881 ( .A(pos_disp_tx), .B(n180), .Z(n2432) );
  AN2 U1882 ( .A(n291), .B(n25), .Z(n2431) );
  AN2 U1883 ( .A(pos_disp_tx), .B(n205), .Z(n2430) );
  AN2 U1884 ( .A(pos_disp_tx), .B(n29), .Z(n2429) );
  AN2 U1885 ( .A(n291), .B(n218), .Z(n2428) );
  AN2 U1886 ( .A(n291), .B(n267), .Z(n2427) );
  AN2 U1887 ( .A(n291), .B(n133), .Z(n2426) );
  AN2 U1888 ( .A(n291), .B(n181), .Z(n2425) );
  AN2 U1889 ( .A(pos_disp_tx), .B(n60), .Z(n2424) );
  AN2 U1890 ( .A(n291), .B(n231), .Z(n2423) );
  AN2 U1891 ( .A(n291), .B(n97), .Z(n2422) );
  AN2 U1892 ( .A(n291), .B(n48), .Z(n2421) );
  AN2 U1893 ( .A(pos_disp_tx), .B(n206), .Z(n2420) );
  AN2 U1894 ( .A(pos_disp_tx), .B(n72), .Z(n2419) );
  AN2 U1895 ( .A(pos_disp_tx), .B(n182), .Z(n2418) );
  AN2 U1896 ( .A(n291), .B(n61), .Z(n2417) );
  AN2 U1897 ( .A(pos_disp_tx), .B(n207), .Z(n2416) );
  AN2 U1898 ( .A(pos_disp_tx), .B(n73), .Z(n2415) );
  AN2 U1899 ( .A(n291), .B(n220), .Z(n2414) );
  AN2 U1900 ( .A(n291), .B(n269), .Z(n2413) );
  AN2 U1901 ( .A(n291), .B(n135), .Z(n2412) );
  AN2 U1902 ( .A(n291), .B(n183), .Z(n2411) );
  AN2 U1903 ( .A(pos_disp_tx), .B(n62), .Z(n2410) );
  AN2 U1904 ( .A(n291), .B(n233), .Z(n2409) );
  AN2 U1905 ( .A(n291), .B(n99), .Z(n2408) );
  AN2 U1906 ( .A(n291), .B(n50), .Z(n2407) );
  AN2 U1907 ( .A(pos_disp_tx), .B(n208), .Z(n2406) );
  AN2 U1908 ( .A(pos_disp_tx), .B(n74), .Z(n2405) );
  AN2 U1909 ( .A(pos_disp_tx), .B(n184), .Z(n2404) );
  AN2 U1910 ( .A(n291), .B(n63), .Z(n2403) );
  AN2 U1911 ( .A(pos_disp_tx), .B(n209), .Z(n2402) );
  AN2 U1912 ( .A(pos_disp_tx), .B(n75), .Z(n2401) );
  AN2 U1913 ( .A(n291), .B(n222), .Z(n2400) );
  AN2 U1914 ( .A(n291), .B(n271), .Z(n2399) );
  AN2 U1915 ( .A(n291), .B(n137), .Z(n2398) );
  AN2 U1916 ( .A(n291), .B(n185), .Z(n2397) );
  AN2 U1917 ( .A(pos_disp_tx), .B(n64), .Z(n2396) );
  AN2 U1918 ( .A(n291), .B(n235), .Z(n2395) );
  AN2 U1919 ( .A(n291), .B(n101), .Z(n2394) );
  AN2 U1920 ( .A(n291), .B(n52), .Z(n2393) );
  AN2 U1921 ( .A(pos_disp_tx), .B(n210), .Z(n2392) );
  AN2 U1922 ( .A(pos_disp_tx), .B(n76), .Z(n2391) );
  AN2 U1923 ( .A(pos_disp_tx), .B(n186), .Z(n2390) );
  AN2 U1924 ( .A(n291), .B(n65), .Z(n2389) );
  AN2 U1925 ( .A(pos_disp_tx), .B(n211), .Z(n2388) );
  AN2 U1926 ( .A(pos_disp_tx), .B(n77), .Z(n2387) );
  AN2 U1927 ( .A(n291), .B(n224), .Z(n2386) );
  AN2 U1928 ( .A(n291), .B(n273), .Z(n2385) );
  AN2 U1929 ( .A(n291), .B(n139), .Z(n2384) );
  AN2 U1930 ( .A(n291), .B(n187), .Z(n2383) );
  AN2 U1931 ( .A(pos_disp_tx), .B(n66), .Z(n2382) );
  AN2 U1932 ( .A(n291), .B(n237), .Z(n2381) );
  AN2 U1933 ( .A(n291), .B(n103), .Z(n2380) );
  AN2 U1934 ( .A(n291), .B(n54), .Z(n2379) );
  AN2 U1935 ( .A(pos_disp_tx), .B(n212), .Z(n2378) );
  AN2 U1936 ( .A(pos_disp_tx), .B(n78), .Z(n2377) );
  AN2 U1937 ( .A(pos_disp_tx), .B(n188), .Z(n2376) );
  AN2 U1938 ( .A(n291), .B(n67), .Z(n2375) );
  AN2 U1939 ( .A(pos_disp_tx), .B(n213), .Z(n2374) );
  AN2 U1940 ( .A(pos_disp_tx), .B(n79), .Z(n2373) );
  AN2 U1941 ( .A(n291), .B(n226), .Z(n2372) );
  AN2 U1942 ( .A(n291), .B(n275), .Z(n2371) );
  AN2 U1943 ( .A(n291), .B(n141), .Z(n2370) );
  AN2 U1944 ( .A(n291), .B(n189), .Z(n2369) );
  AN2 U1945 ( .A(pos_disp_tx), .B(n68), .Z(n2368) );
  AN2 U1946 ( .A(n291), .B(n239), .Z(n2367) );
  AN2 U1947 ( .A(n291), .B(n105), .Z(n2366) );
  AN2 U1948 ( .A(n291), .B(n56), .Z(n2365) );
  AN2 U1949 ( .A(pos_disp_tx), .B(n214), .Z(n2364) );
  AN2 U1950 ( .A(pos_disp_tx), .B(n80), .Z(n2363) );
  AN2 U1951 ( .A(pos_disp_tx), .B(n190), .Z(n2362) );
  AN2 U1952 ( .A(n291), .B(n69), .Z(n2361) );
  AN2 U1953 ( .A(pos_disp_tx), .B(n215), .Z(n2360) );
  AN2 U1954 ( .A(pos_disp_tx), .B(n81), .Z(n2359) );
  AN2 U1955 ( .A(n291), .B(n228), .Z(n2358) );
  AN2 U1956 ( .A(n291), .B(n277), .Z(n2357) );
  AN2 U1957 ( .A(n291), .B(n143), .Z(n2356) );
  AN2 U1958 ( .A(n291), .B(n191), .Z(n2355) );
  AN2 U1959 ( .A(pos_disp_tx), .B(n70), .Z(n2354) );
  AN2 U1960 ( .A(n291), .B(n241), .Z(n2353) );
  AN2 U1961 ( .A(n291), .B(n107), .Z(n2352) );
  AN2 U1962 ( .A(n291), .B(n58), .Z(n2351) );
  AN2 U1963 ( .A(pos_disp_tx), .B(n216), .Z(n2350) );
  AN2 U1964 ( .A(pos_disp_tx), .B(n82), .Z(n2349) );
  AN2 U1965 ( .A(pos_disp_tx), .B(n192), .Z(n2348) );
  AN2 U1966 ( .A(n291), .B(n71), .Z(n2347) );
  AN2 U1967 ( .A(pos_disp_tx), .B(n217), .Z(n2346) );
  AN2 U1968 ( .A(pos_disp_tx), .B(n83), .Z(n2345) );
  AN2 U1969 ( .A(n291), .B(n230), .Z(n2344) );
  AN2 U1970 ( .A(n291), .B(n279), .Z(n2343) );
  AN2 U1971 ( .A(n291), .B(n145), .Z(n2342) );
  AN2 U1972 ( .A(n291), .B(N239), .Z(n2341) );
  OR2 U1973 ( .A(n2339), .B(n2340), .Z(N837) );
  OR2 U1974 ( .A(n2337), .B(n2338), .Z(n2340) );
  OR2 U1975 ( .A(n2335), .B(n2336), .Z(n2339) );
  OR2 U1976 ( .A(n2334), .B(n2285), .Z(n2338) );
  OR2 U1977 ( .A(n2332), .B(n2333), .Z(n2337) );
  OR2 U1978 ( .A(n2330), .B(n2331), .Z(n2336) );
  OR2 U1979 ( .A(n2328), .B(n2329), .Z(n2335) );
  OR2 U1980 ( .A(n2326), .B(n2327), .Z(n2334) );
  OR2 U1981 ( .A(n2324), .B(n2325), .Z(n2333) );
  OR2 U1982 ( .A(n2322), .B(n2323), .Z(n2332) );
  OR2 U1983 ( .A(n2320), .B(n2321), .Z(n2331) );
  OR2 U1984 ( .A(n2318), .B(n2319), .Z(n2330) );
  OR2 U1985 ( .A(n2316), .B(n2317), .Z(n2329) );
  OR2 U1986 ( .A(n2314), .B(n2315), .Z(n2328) );
  OR2 U1987 ( .A(n2312), .B(n2313), .Z(n2327) );
  OR2 U1988 ( .A(n2310), .B(n2311), .Z(n2326) );
  OR2 U1989 ( .A(n2308), .B(n2309), .Z(n2325) );
  OR2 U1990 ( .A(n2306), .B(n2307), .Z(n2324) );
  OR2 U1991 ( .A(n2304), .B(n2305), .Z(n2323) );
  OR2 U1992 ( .A(n2302), .B(n2303), .Z(n2322) );
  OR2 U1993 ( .A(n2300), .B(n2301), .Z(n2321) );
  OR2 U1994 ( .A(n2298), .B(n2299), .Z(n2320) );
  OR2 U1995 ( .A(n2296), .B(n2297), .Z(n2319) );
  OR2 U1996 ( .A(n2294), .B(n2295), .Z(n2318) );
  OR2 U1997 ( .A(n2292), .B(n2293), .Z(n2317) );
  OR2 U1998 ( .A(n2290), .B(n2291), .Z(n2316) );
  OR2 U1999 ( .A(n2288), .B(n2289), .Z(n2315) );
  OR2 U2000 ( .A(n2286), .B(n2287), .Z(n2314) );
  OR2 U2001 ( .A(n2283), .B(n2284), .Z(n2313) );
  OR2 U2002 ( .A(n2281), .B(n2282), .Z(n2312) );
  OR2 U2003 ( .A(n2279), .B(n2280), .Z(n2311) );
  OR2 U2004 ( .A(n2277), .B(n2278), .Z(n2310) );
  OR2 U2005 ( .A(n2275), .B(n2276), .Z(n2309) );
  OR2 U2006 ( .A(n2273), .B(n2274), .Z(n2308) );
  OR2 U2007 ( .A(n2271), .B(n2272), .Z(n2307) );
  OR2 U2008 ( .A(n2269), .B(n2270), .Z(n2306) );
  OR2 U2009 ( .A(n2267), .B(n2268), .Z(n2305) );
  OR2 U2010 ( .A(n2265), .B(n2266), .Z(n2304) );
  OR2 U2011 ( .A(n2263), .B(n2264), .Z(n2303) );
  OR2 U2012 ( .A(n2261), .B(n2262), .Z(n2302) );
  OR2 U2013 ( .A(n2259), .B(n2260), .Z(n2301) );
  OR2 U2014 ( .A(n2257), .B(n2258), .Z(n2300) );
  OR2 U2015 ( .A(n2255), .B(n2256), .Z(n2299) );
  OR2 U2016 ( .A(n2253), .B(n2254), .Z(n2298) );
  OR2 U2017 ( .A(n2251), .B(n2252), .Z(n2297) );
  OR2 U2018 ( .A(n2249), .B(n2250), .Z(n2296) );
  OR2 U2019 ( .A(n2247), .B(n2248), .Z(n2295) );
  OR2 U2020 ( .A(n2245), .B(n2246), .Z(n2294) );
  OR2 U2021 ( .A(n2243), .B(n2244), .Z(n2293) );
  OR2 U2022 ( .A(n2241), .B(n2242), .Z(n2292) );
  OR2 U2023 ( .A(n2239), .B(n2240), .Z(n2291) );
  OR2 U2024 ( .A(n2237), .B(n2238), .Z(n2290) );
  OR2 U2025 ( .A(n2235), .B(n2236), .Z(n2289) );
  OR2 U2026 ( .A(n2233), .B(n2234), .Z(n2288) );
  OR2 U2027 ( .A(n2231), .B(n2232), .Z(n2287) );
  OR2 U2028 ( .A(n2230), .B(n2120), .Z(n2286) );
  OR2 U2029 ( .A(n2228), .B(n2229), .Z(n2285) );
  OR2 U2030 ( .A(n2226), .B(n2227), .Z(n2284) );
  OR2 U2031 ( .A(n2224), .B(n2225), .Z(n2283) );
  OR2 U2032 ( .A(n2222), .B(n2223), .Z(n2282) );
  OR2 U2033 ( .A(n2220), .B(n2221), .Z(n2281) );
  OR2 U2034 ( .A(n2218), .B(n2219), .Z(n2280) );
  OR2 U2035 ( .A(n2216), .B(n2217), .Z(n2279) );
  OR2 U2036 ( .A(n2214), .B(n2215), .Z(n2278) );
  OR2 U2037 ( .A(n2212), .B(n2213), .Z(n2277) );
  OR2 U2038 ( .A(n2210), .B(n2211), .Z(n2276) );
  OR2 U2039 ( .A(n2208), .B(n2209), .Z(n2275) );
  OR2 U2040 ( .A(n2206), .B(n2207), .Z(n2274) );
  OR2 U2041 ( .A(n2204), .B(n2205), .Z(n2273) );
  OR2 U2042 ( .A(n2202), .B(n2203), .Z(n2272) );
  OR2 U2043 ( .A(n2200), .B(n2201), .Z(n2271) );
  OR2 U2044 ( .A(n2198), .B(n2199), .Z(n2270) );
  OR2 U2045 ( .A(n2196), .B(n2197), .Z(n2269) );
  OR2 U2046 ( .A(n2194), .B(n2195), .Z(n2268) );
  OR2 U2047 ( .A(n2192), .B(n2193), .Z(n2267) );
  OR2 U2048 ( .A(n2190), .B(n2191), .Z(n2266) );
  OR2 U2049 ( .A(n2188), .B(n2189), .Z(n2265) );
  OR2 U2050 ( .A(n2186), .B(n2187), .Z(n2264) );
  OR2 U2051 ( .A(n2184), .B(n2185), .Z(n2263) );
  OR2 U2052 ( .A(n2182), .B(n2183), .Z(n2262) );
  OR2 U2053 ( .A(n2180), .B(n2181), .Z(n2261) );
  OR2 U2054 ( .A(n2178), .B(n2179), .Z(n2260) );
  OR2 U2055 ( .A(n2176), .B(n2177), .Z(n2259) );
  OR2 U2056 ( .A(n2174), .B(n2175), .Z(n2258) );
  OR2 U2057 ( .A(n2172), .B(n2173), .Z(n2257) );
  OR2 U2058 ( .A(n2170), .B(n2171), .Z(n2256) );
  OR2 U2059 ( .A(n2168), .B(n2169), .Z(n2255) );
  OR2 U2060 ( .A(n2166), .B(n2167), .Z(n2254) );
  OR2 U2061 ( .A(n2164), .B(n2165), .Z(n2253) );
  OR2 U2062 ( .A(n2162), .B(n2163), .Z(n2252) );
  OR2 U2063 ( .A(n2160), .B(n2161), .Z(n2251) );
  OR2 U2064 ( .A(n2158), .B(n2159), .Z(n2250) );
  OR2 U2065 ( .A(n2156), .B(n2157), .Z(n2249) );
  OR2 U2066 ( .A(n2154), .B(n2155), .Z(n2248) );
  OR2 U2067 ( .A(n2152), .B(n2153), .Z(n2247) );
  OR2 U2068 ( .A(n2150), .B(n2151), .Z(n2246) );
  OR2 U2069 ( .A(n2148), .B(n2149), .Z(n2245) );
  OR2 U2070 ( .A(n2146), .B(n2147), .Z(n2244) );
  OR2 U2071 ( .A(n2144), .B(n2145), .Z(n2243) );
  OR2 U2072 ( .A(n2142), .B(n2143), .Z(n2242) );
  OR2 U2073 ( .A(n2140), .B(n2141), .Z(n2241) );
  OR2 U2074 ( .A(n2138), .B(n2139), .Z(n2240) );
  OR2 U2075 ( .A(n2136), .B(n2137), .Z(n2239) );
  OR2 U2076 ( .A(n2134), .B(n2135), .Z(n2238) );
  OR2 U2077 ( .A(n2132), .B(n2133), .Z(n2237) );
  OR2 U2078 ( .A(n2130), .B(n2131), .Z(n2236) );
  OR2 U2079 ( .A(n2128), .B(n2129), .Z(n2235) );
  OR2 U2080 ( .A(n2126), .B(n2127), .Z(n2234) );
  OR2 U2081 ( .A(n2125), .B(N1027), .Z(n2233) );
  OR2 U2082 ( .A(n2123), .B(n2124), .Z(n2232) );
  OR2 U2083 ( .A(n2121), .B(n2122), .Z(n2231) );
  OR2 U2084 ( .A(n2118), .B(n2119), .Z(n2230) );
  AN2 U2085 ( .A(n291), .B(N8311), .Z(n2229) );
  AN2 U2086 ( .A(n291), .B(n153), .Z(n2228) );
  AN2 U2087 ( .A(n291), .B(n33), .Z(n2227) );
  AN2 U2088 ( .A(n291), .B(n19), .Z(n2226) );
  AN2 U2089 ( .A(n291), .B(n172), .Z(n2225) );
  AN2 U2090 ( .A(n291), .B(n26), .Z(n2224) );
  AN2 U2091 ( .A(n291), .B(n178), .Z(n2223) );
  AN2 U2092 ( .A(n291), .B(n23), .Z(n2222) );
  AN2 U2093 ( .A(pos_disp_tx), .B(n173), .Z(n2221) );
  AN2 U2094 ( .A(pos_disp_tx), .B(n27), .Z(n2220) );
  AN2 U2095 ( .A(pos_disp_tx), .B(n176), .Z(n2219) );
  AN2 U2096 ( .A(pos_disp_tx), .B(n166), .Z(n2218) );
  AN2 U2097 ( .A(pos_disp_tx), .B(n44), .Z(n2217) );
  AN2 U2098 ( .A(n291), .B(n179), .Z(n2216) );
  AN2 U2099 ( .A(n291), .B(n24), .Z(n2215) );
  AN2 U2100 ( .A(n291), .B(n155), .Z(n2214) );
  AN2 U2101 ( .A(n291), .B(n35), .Z(n2213) );
  AN2 U2102 ( .A(n291), .B(n21), .Z(n2212) );
  AN2 U2103 ( .A(n291), .B(n174), .Z(n2211) );
  AN2 U2104 ( .A(n291), .B(n28), .Z(n2210) );
  AN2 U2105 ( .A(n291), .B(n180), .Z(n2209) );
  AN2 U2106 ( .A(n291), .B(n25), .Z(n2208) );
  AN2 U2107 ( .A(pos_disp_tx), .B(n205), .Z(n2207) );
  AN2 U2108 ( .A(pos_disp_tx), .B(n29), .Z(n2206) );
  AN2 U2109 ( .A(pos_disp_tx), .B(n218), .Z(n2205) );
  AN2 U2110 ( .A(pos_disp_tx), .B(n267), .Z(n2204) );
  AN2 U2111 ( .A(pos_disp_tx), .B(n133), .Z(n2203) );
  AN2 U2112 ( .A(n291), .B(n181), .Z(n2202) );
  AN2 U2113 ( .A(n291), .B(n60), .Z(n2201) );
  AN2 U2114 ( .A(n291), .B(n231), .Z(n2200) );
  AN2 U2115 ( .A(n291), .B(n97), .Z(n2199) );
  AN2 U2116 ( .A(n291), .B(n48), .Z(n2198) );
  AN2 U2117 ( .A(n291), .B(n206), .Z(n2197) );
  AN2 U2118 ( .A(n291), .B(n72), .Z(n2196) );
  AN2 U2119 ( .A(n291), .B(n182), .Z(n2195) );
  AN2 U2120 ( .A(n291), .B(n61), .Z(n2194) );
  AN2 U2121 ( .A(pos_disp_tx), .B(n207), .Z(n2193) );
  AN2 U2122 ( .A(pos_disp_tx), .B(n73), .Z(n2192) );
  AN2 U2123 ( .A(pos_disp_tx), .B(n220), .Z(n2191) );
  AN2 U2124 ( .A(pos_disp_tx), .B(n269), .Z(n2190) );
  AN2 U2125 ( .A(pos_disp_tx), .B(n135), .Z(n2189) );
  AN2 U2126 ( .A(n291), .B(n183), .Z(n2188) );
  AN2 U2127 ( .A(n291), .B(n62), .Z(n2187) );
  AN2 U2128 ( .A(n291), .B(n233), .Z(n2186) );
  AN2 U2129 ( .A(n291), .B(n99), .Z(n2185) );
  AN2 U2130 ( .A(n291), .B(n50), .Z(n2184) );
  AN2 U2131 ( .A(n291), .B(n208), .Z(n2183) );
  AN2 U2132 ( .A(n291), .B(n74), .Z(n2182) );
  AN2 U2133 ( .A(n291), .B(n184), .Z(n2181) );
  AN2 U2134 ( .A(n291), .B(n63), .Z(n2180) );
  AN2 U2135 ( .A(pos_disp_tx), .B(n209), .Z(n2179) );
  AN2 U2136 ( .A(pos_disp_tx), .B(n75), .Z(n2178) );
  AN2 U2137 ( .A(pos_disp_tx), .B(n222), .Z(n2177) );
  AN2 U2138 ( .A(pos_disp_tx), .B(n271), .Z(n2176) );
  AN2 U2139 ( .A(pos_disp_tx), .B(n137), .Z(n2175) );
  AN2 U2140 ( .A(n291), .B(n185), .Z(n2174) );
  AN2 U2141 ( .A(n291), .B(n64), .Z(n2173) );
  AN2 U2142 ( .A(n291), .B(n235), .Z(n2172) );
  AN2 U2143 ( .A(n291), .B(n101), .Z(n2171) );
  AN2 U2144 ( .A(n291), .B(n52), .Z(n2170) );
  AN2 U2145 ( .A(n291), .B(n210), .Z(n2169) );
  AN2 U2146 ( .A(n291), .B(n76), .Z(n2168) );
  AN2 U2147 ( .A(n291), .B(n186), .Z(n2167) );
  AN2 U2148 ( .A(n291), .B(n65), .Z(n2166) );
  AN2 U2149 ( .A(pos_disp_tx), .B(n211), .Z(n2165) );
  AN2 U2150 ( .A(pos_disp_tx), .B(n77), .Z(n2164) );
  AN2 U2151 ( .A(pos_disp_tx), .B(n224), .Z(n2163) );
  AN2 U2152 ( .A(pos_disp_tx), .B(n273), .Z(n2162) );
  AN2 U2153 ( .A(pos_disp_tx), .B(n139), .Z(n2161) );
  AN2 U2154 ( .A(n291), .B(n187), .Z(n2160) );
  AN2 U2155 ( .A(n291), .B(n66), .Z(n2159) );
  AN2 U2156 ( .A(n291), .B(n237), .Z(n2158) );
  AN2 U2157 ( .A(n291), .B(n103), .Z(n2157) );
  AN2 U2158 ( .A(n291), .B(n54), .Z(n2156) );
  AN2 U2159 ( .A(n291), .B(n212), .Z(n2155) );
  AN2 U2160 ( .A(n291), .B(n78), .Z(n2154) );
  AN2 U2161 ( .A(n291), .B(n188), .Z(n2153) );
  AN2 U2162 ( .A(n291), .B(n67), .Z(n2152) );
  AN2 U2163 ( .A(pos_disp_tx), .B(n213), .Z(n2151) );
  AN2 U2164 ( .A(pos_disp_tx), .B(n79), .Z(n2150) );
  AN2 U2165 ( .A(pos_disp_tx), .B(n226), .Z(n2149) );
  AN2 U2166 ( .A(pos_disp_tx), .B(n275), .Z(n2148) );
  AN2 U2167 ( .A(pos_disp_tx), .B(n141), .Z(n2147) );
  AN2 U2168 ( .A(n291), .B(n189), .Z(n2146) );
  AN2 U2169 ( .A(n291), .B(n68), .Z(n2145) );
  AN2 U2170 ( .A(n291), .B(n239), .Z(n2144) );
  AN2 U2171 ( .A(n291), .B(n105), .Z(n2143) );
  AN2 U2172 ( .A(n291), .B(n56), .Z(n2142) );
  AN2 U2173 ( .A(n291), .B(n214), .Z(n2141) );
  AN2 U2174 ( .A(n291), .B(n80), .Z(n2140) );
  AN2 U2175 ( .A(n291), .B(n190), .Z(n2139) );
  AN2 U2176 ( .A(n291), .B(n69), .Z(n2138) );
  AN2 U2177 ( .A(pos_disp_tx), .B(n215), .Z(n2137) );
  AN2 U2178 ( .A(pos_disp_tx), .B(n81), .Z(n2136) );
  AN2 U2179 ( .A(pos_disp_tx), .B(n228), .Z(n2135) );
  AN2 U2180 ( .A(pos_disp_tx), .B(n277), .Z(n2134) );
  AN2 U2181 ( .A(pos_disp_tx), .B(n143), .Z(n2133) );
  AN2 U2182 ( .A(n291), .B(n191), .Z(n2132) );
  AN2 U2183 ( .A(n291), .B(n70), .Z(n2131) );
  AN2 U2184 ( .A(n291), .B(n241), .Z(n2130) );
  AN2 U2185 ( .A(n291), .B(n107), .Z(n2129) );
  AN2 U2186 ( .A(n291), .B(n58), .Z(n2128) );
  AN2 U2187 ( .A(n291), .B(n216), .Z(n2127) );
  AN2 U2188 ( .A(n291), .B(n82), .Z(n2126) );
  AN2 U2189 ( .A(n291), .B(n192), .Z(n2125) );
  AN2 U2190 ( .A(n291), .B(n71), .Z(n2124) );
  AN2 U2191 ( .A(pos_disp_tx), .B(n217), .Z(n2123) );
  AN2 U2192 ( .A(pos_disp_tx), .B(n83), .Z(n2122) );
  AN2 U2193 ( .A(pos_disp_tx), .B(n230), .Z(n2121) );
  AN2 U2194 ( .A(pos_disp_tx), .B(n279), .Z(n2120) );
  AN2 U2195 ( .A(pos_disp_tx), .B(n145), .Z(n2119) );
  AN2 U2196 ( .A(n291), .B(N239), .Z(n2118) );
  OR2 U2197 ( .A(n2116), .B(n2117), .Z(N836) );
  OR2 U2198 ( .A(n2114), .B(n2115), .Z(n2117) );
  OR2 U2199 ( .A(n2112), .B(n2113), .Z(n2116) );
  OR2 U2200 ( .A(n2111), .B(n2062), .Z(n2115) );
  OR2 U2201 ( .A(n2109), .B(n2110), .Z(n2114) );
  OR2 U2202 ( .A(n2107), .B(n2108), .Z(n2113) );
  OR2 U2203 ( .A(n2105), .B(n2106), .Z(n2112) );
  OR2 U2204 ( .A(n2103), .B(n2104), .Z(n2111) );
  OR2 U2205 ( .A(n2101), .B(n2102), .Z(n2110) );
  OR2 U2206 ( .A(n2099), .B(n2100), .Z(n2109) );
  OR2 U2207 ( .A(n2097), .B(n2098), .Z(n2108) );
  OR2 U2208 ( .A(n2095), .B(n2096), .Z(n2107) );
  OR2 U2209 ( .A(n2093), .B(n2094), .Z(n2106) );
  OR2 U2210 ( .A(n2091), .B(n2092), .Z(n2105) );
  OR2 U2211 ( .A(n2089), .B(n2090), .Z(n2104) );
  OR2 U2212 ( .A(n2087), .B(n2088), .Z(n2103) );
  OR2 U2213 ( .A(n2085), .B(n2086), .Z(n2102) );
  OR2 U2214 ( .A(n2083), .B(n2084), .Z(n2101) );
  OR2 U2215 ( .A(n2081), .B(n2082), .Z(n2100) );
  OR2 U2216 ( .A(n2079), .B(n2080), .Z(n2099) );
  OR2 U2217 ( .A(n2077), .B(n2078), .Z(n2098) );
  OR2 U2218 ( .A(n2075), .B(n2076), .Z(n2097) );
  OR2 U2219 ( .A(n2073), .B(n2074), .Z(n2096) );
  OR2 U2220 ( .A(n2071), .B(n2072), .Z(n2095) );
  OR2 U2221 ( .A(n2069), .B(n2070), .Z(n2094) );
  OR2 U2222 ( .A(n2067), .B(n2068), .Z(n2093) );
  OR2 U2223 ( .A(n2065), .B(n2066), .Z(n2092) );
  OR2 U2224 ( .A(n2063), .B(n2064), .Z(n2091) );
  OR2 U2225 ( .A(n2060), .B(n2061), .Z(n2090) );
  OR2 U2226 ( .A(n2058), .B(n2059), .Z(n2089) );
  OR2 U2227 ( .A(n2056), .B(n2057), .Z(n2088) );
  OR2 U2228 ( .A(n2054), .B(n2055), .Z(n2087) );
  OR2 U2229 ( .A(n2052), .B(n2053), .Z(n2086) );
  OR2 U2230 ( .A(n2050), .B(n2051), .Z(n2085) );
  OR2 U2231 ( .A(n2048), .B(n2049), .Z(n2084) );
  OR2 U2232 ( .A(n2046), .B(n2047), .Z(n2083) );
  OR2 U2233 ( .A(n2044), .B(n2045), .Z(n2082) );
  OR2 U2234 ( .A(n2042), .B(n2043), .Z(n2081) );
  OR2 U2235 ( .A(n2040), .B(n2041), .Z(n2080) );
  OR2 U2236 ( .A(n2038), .B(n2039), .Z(n2079) );
  OR2 U2237 ( .A(n2036), .B(n2037), .Z(n2078) );
  OR2 U2238 ( .A(n2034), .B(n2035), .Z(n2077) );
  OR2 U2239 ( .A(n2032), .B(n2033), .Z(n2076) );
  OR2 U2240 ( .A(n2030), .B(n2031), .Z(n2075) );
  OR2 U2241 ( .A(n2028), .B(n2029), .Z(n2074) );
  OR2 U2242 ( .A(n2026), .B(n2027), .Z(n2073) );
  OR2 U2243 ( .A(n2024), .B(n2025), .Z(n2072) );
  OR2 U2244 ( .A(n2022), .B(n2023), .Z(n2071) );
  OR2 U2245 ( .A(n2020), .B(n2021), .Z(n2070) );
  OR2 U2246 ( .A(n2018), .B(n2019), .Z(n2069) );
  OR2 U2247 ( .A(n2016), .B(n2017), .Z(n2068) );
  OR2 U2248 ( .A(n2014), .B(n2015), .Z(n2067) );
  OR2 U2249 ( .A(n2012), .B(n2013), .Z(n2066) );
  OR2 U2250 ( .A(n2010), .B(n2011), .Z(n2065) );
  OR2 U2251 ( .A(n2009), .B(n1900), .Z(n2064) );
  OR2 U2252 ( .A(n2007), .B(n2008), .Z(n2063) );
  OR2 U2253 ( .A(n2005), .B(n2006), .Z(n2062) );
  OR2 U2254 ( .A(n2003), .B(n2004), .Z(n2061) );
  OR2 U2255 ( .A(n2001), .B(n2002), .Z(n2060) );
  OR2 U2256 ( .A(n1999), .B(n2000), .Z(n2059) );
  OR2 U2257 ( .A(n1997), .B(n1998), .Z(n2058) );
  OR2 U2258 ( .A(n1995), .B(n1996), .Z(n2057) );
  OR2 U2259 ( .A(n1993), .B(n1994), .Z(n2056) );
  OR2 U2260 ( .A(n1991), .B(n1992), .Z(n2055) );
  OR2 U2261 ( .A(n1989), .B(n1990), .Z(n2054) );
  OR2 U2262 ( .A(n1987), .B(n1988), .Z(n2053) );
  OR2 U2263 ( .A(n1985), .B(n1986), .Z(n2052) );
  OR2 U2264 ( .A(n1983), .B(n1984), .Z(n2051) );
  OR2 U2265 ( .A(n1981), .B(n1982), .Z(n2050) );
  OR2 U2266 ( .A(n1979), .B(n1980), .Z(n2049) );
  OR2 U2267 ( .A(n1977), .B(n1978), .Z(n2048) );
  OR2 U2268 ( .A(n1975), .B(n1976), .Z(n2047) );
  OR2 U2269 ( .A(n1973), .B(n1974), .Z(n2046) );
  OR2 U2270 ( .A(n1971), .B(n1972), .Z(n2045) );
  OR2 U2271 ( .A(n1969), .B(n1970), .Z(n2044) );
  OR2 U2272 ( .A(n1967), .B(n1968), .Z(n2043) );
  OR2 U2273 ( .A(n1965), .B(n1966), .Z(n2042) );
  OR2 U2274 ( .A(n1963), .B(n1964), .Z(n2041) );
  OR2 U2275 ( .A(n1961), .B(n1962), .Z(n2040) );
  OR2 U2276 ( .A(n1959), .B(n1960), .Z(n2039) );
  OR2 U2277 ( .A(n1957), .B(n1958), .Z(n2038) );
  OR2 U2278 ( .A(n1955), .B(n1956), .Z(n2037) );
  OR2 U2279 ( .A(n1953), .B(n1954), .Z(n2036) );
  OR2 U2280 ( .A(n1951), .B(n1952), .Z(n2035) );
  OR2 U2281 ( .A(n1949), .B(n1950), .Z(n2034) );
  OR2 U2282 ( .A(n1947), .B(n1948), .Z(n2033) );
  OR2 U2283 ( .A(n1945), .B(n1946), .Z(n2032) );
  OR2 U2284 ( .A(n1943), .B(n1944), .Z(n2031) );
  OR2 U2285 ( .A(n1941), .B(n1942), .Z(n2030) );
  OR2 U2286 ( .A(n1939), .B(n1940), .Z(n2029) );
  OR2 U2287 ( .A(n1937), .B(n1938), .Z(n2028) );
  OR2 U2288 ( .A(n1935), .B(n1936), .Z(n2027) );
  OR2 U2289 ( .A(n1933), .B(n1934), .Z(n2026) );
  OR2 U2290 ( .A(n1931), .B(n1932), .Z(n2025) );
  OR2 U2291 ( .A(n1929), .B(n1930), .Z(n2024) );
  OR2 U2292 ( .A(n1927), .B(n1928), .Z(n2023) );
  OR2 U2293 ( .A(n1925), .B(n1926), .Z(n2022) );
  OR2 U2294 ( .A(n1923), .B(n1924), .Z(n2021) );
  OR2 U2295 ( .A(n1921), .B(n1922), .Z(n2020) );
  OR2 U2296 ( .A(n1919), .B(n1920), .Z(n2019) );
  OR2 U2297 ( .A(n1917), .B(n1918), .Z(n2018) );
  OR2 U2298 ( .A(n1915), .B(n1916), .Z(n2017) );
  OR2 U2299 ( .A(n1913), .B(n1914), .Z(n2016) );
  OR2 U2300 ( .A(n1911), .B(n1912), .Z(n2015) );
  OR2 U2301 ( .A(n1909), .B(n1910), .Z(n2014) );
  OR2 U2302 ( .A(n1907), .B(n1908), .Z(n2013) );
  OR2 U2303 ( .A(n1905), .B(n1906), .Z(n2012) );
  OR2 U2304 ( .A(n1903), .B(n1904), .Z(n2011) );
  OR2 U2305 ( .A(n1901), .B(n1902), .Z(n2010) );
  OR2 U2306 ( .A(n1898), .B(n1899), .Z(n2009) );
  OR2 U2307 ( .A(n1897), .B(N976), .Z(n2008) );
  OR2 U2308 ( .A(n1895), .B(n1896), .Z(n2007) );
  AN2 U2309 ( .A(n291), .B(N8311), .Z(n2006) );
  AN2 U2310 ( .A(pos_disp_tx), .B(n153), .Z(n2005) );
  AN2 U2311 ( .A(pos_disp_tx), .B(n33), .Z(n2004) );
  AN2 U2312 ( .A(pos_disp_tx), .B(n19), .Z(n2003) );
  AN2 U2313 ( .A(n291), .B(n172), .Z(n2002) );
  AN2 U2314 ( .A(pos_disp_tx), .B(n26), .Z(n2001) );
  AN2 U2315 ( .A(n291), .B(n178), .Z(n2000) );
  AN2 U2316 ( .A(n291), .B(n23), .Z(n1999) );
  AN2 U2317 ( .A(n291), .B(n173), .Z(n1998) );
  AN2 U2318 ( .A(pos_disp_tx), .B(n27), .Z(n1997) );
  AN2 U2319 ( .A(n291), .B(n176), .Z(n1996) );
  AN2 U2320 ( .A(n291), .B(n166), .Z(n1995) );
  AN2 U2321 ( .A(n291), .B(n44), .Z(n1994) );
  AN2 U2322 ( .A(n291), .B(n179), .Z(n1993) );
  AN2 U2323 ( .A(n291), .B(n24), .Z(n1992) );
  AN2 U2324 ( .A(pos_disp_tx), .B(n155), .Z(n1991) );
  AN2 U2325 ( .A(pos_disp_tx), .B(n35), .Z(n1990) );
  AN2 U2326 ( .A(pos_disp_tx), .B(n21), .Z(n1989) );
  AN2 U2327 ( .A(n291), .B(n174), .Z(n1988) );
  AN2 U2328 ( .A(pos_disp_tx), .B(n28), .Z(n1987) );
  AN2 U2329 ( .A(n291), .B(n180), .Z(n1986) );
  AN2 U2330 ( .A(n291), .B(n25), .Z(n1985) );
  AN2 U2331 ( .A(n291), .B(n205), .Z(n1984) );
  AN2 U2332 ( .A(pos_disp_tx), .B(n29), .Z(n1983) );
  AN2 U2333 ( .A(n291), .B(n218), .Z(n1982) );
  AN2 U2334 ( .A(n291), .B(n267), .Z(n1981) );
  AN2 U2335 ( .A(n291), .B(n133), .Z(n1980) );
  AN2 U2336 ( .A(n291), .B(n181), .Z(n1979) );
  AN2 U2337 ( .A(n291), .B(n60), .Z(n1978) );
  AN2 U2338 ( .A(pos_disp_tx), .B(n231), .Z(n1977) );
  AN2 U2339 ( .A(pos_disp_tx), .B(n97), .Z(n1976) );
  AN2 U2340 ( .A(pos_disp_tx), .B(n48), .Z(n1975) );
  AN2 U2341 ( .A(n291), .B(n206), .Z(n1974) );
  AN2 U2342 ( .A(pos_disp_tx), .B(n72), .Z(n1973) );
  AN2 U2343 ( .A(n291), .B(n182), .Z(n1972) );
  AN2 U2344 ( .A(n291), .B(n61), .Z(n1971) );
  AN2 U2345 ( .A(n291), .B(n207), .Z(n1970) );
  AN2 U2346 ( .A(pos_disp_tx), .B(n73), .Z(n1969) );
  AN2 U2347 ( .A(n291), .B(n220), .Z(n1968) );
  AN2 U2348 ( .A(n291), .B(n269), .Z(n1967) );
  AN2 U2349 ( .A(n291), .B(n135), .Z(n1966) );
  AN2 U2350 ( .A(n291), .B(n183), .Z(n1965) );
  AN2 U2351 ( .A(n291), .B(n62), .Z(n1964) );
  AN2 U2352 ( .A(pos_disp_tx), .B(n233), .Z(n1963) );
  AN2 U2353 ( .A(pos_disp_tx), .B(n99), .Z(n1962) );
  AN2 U2354 ( .A(pos_disp_tx), .B(n50), .Z(n1961) );
  AN2 U2355 ( .A(n291), .B(n208), .Z(n1960) );
  AN2 U2356 ( .A(pos_disp_tx), .B(n74), .Z(n1959) );
  AN2 U2357 ( .A(n291), .B(n184), .Z(n1958) );
  AN2 U2358 ( .A(n291), .B(n63), .Z(n1957) );
  AN2 U2359 ( .A(n291), .B(n209), .Z(n1956) );
  AN2 U2360 ( .A(pos_disp_tx), .B(n75), .Z(n1955) );
  AN2 U2361 ( .A(n291), .B(n222), .Z(n1954) );
  AN2 U2362 ( .A(n291), .B(n271), .Z(n1953) );
  AN2 U2363 ( .A(n291), .B(n137), .Z(n1952) );
  AN2 U2364 ( .A(n291), .B(n185), .Z(n1951) );
  AN2 U2365 ( .A(n291), .B(n64), .Z(n1950) );
  AN2 U2366 ( .A(pos_disp_tx), .B(n235), .Z(n1949) );
  AN2 U2367 ( .A(pos_disp_tx), .B(n101), .Z(n1948) );
  AN2 U2368 ( .A(pos_disp_tx), .B(n52), .Z(n1947) );
  AN2 U2369 ( .A(n291), .B(n210), .Z(n1946) );
  AN2 U2370 ( .A(pos_disp_tx), .B(n76), .Z(n1945) );
  AN2 U2371 ( .A(n291), .B(n186), .Z(n1944) );
  AN2 U2372 ( .A(n291), .B(n65), .Z(n1943) );
  AN2 U2373 ( .A(n291), .B(n211), .Z(n1942) );
  AN2 U2374 ( .A(pos_disp_tx), .B(n77), .Z(n1941) );
  AN2 U2375 ( .A(n291), .B(n224), .Z(n1940) );
  AN2 U2376 ( .A(n291), .B(n273), .Z(n1939) );
  AN2 U2377 ( .A(n291), .B(n139), .Z(n1938) );
  AN2 U2378 ( .A(n291), .B(n187), .Z(n1937) );
  AN2 U2379 ( .A(n291), .B(n66), .Z(n1936) );
  AN2 U2380 ( .A(pos_disp_tx), .B(n237), .Z(n1935) );
  AN2 U2381 ( .A(pos_disp_tx), .B(n103), .Z(n1934) );
  AN2 U2382 ( .A(pos_disp_tx), .B(n54), .Z(n1933) );
  AN2 U2383 ( .A(n291), .B(n212), .Z(n1932) );
  AN2 U2384 ( .A(pos_disp_tx), .B(n78), .Z(n1931) );
  AN2 U2385 ( .A(n291), .B(n188), .Z(n1930) );
  AN2 U2386 ( .A(n291), .B(n67), .Z(n1929) );
  AN2 U2387 ( .A(n291), .B(n213), .Z(n1928) );
  AN2 U2388 ( .A(pos_disp_tx), .B(n79), .Z(n1927) );
  AN2 U2389 ( .A(n291), .B(n226), .Z(n1926) );
  AN2 U2390 ( .A(n291), .B(n275), .Z(n1925) );
  AN2 U2391 ( .A(n291), .B(n141), .Z(n1924) );
  AN2 U2392 ( .A(n291), .B(n189), .Z(n1923) );
  AN2 U2393 ( .A(n291), .B(n68), .Z(n1922) );
  AN2 U2394 ( .A(pos_disp_tx), .B(n239), .Z(n1921) );
  AN2 U2395 ( .A(pos_disp_tx), .B(n105), .Z(n1920) );
  AN2 U2396 ( .A(pos_disp_tx), .B(n56), .Z(n1919) );
  AN2 U2397 ( .A(n291), .B(n214), .Z(n1918) );
  AN2 U2398 ( .A(pos_disp_tx), .B(n80), .Z(n1917) );
  AN2 U2399 ( .A(n291), .B(n190), .Z(n1916) );
  AN2 U2400 ( .A(n291), .B(n69), .Z(n1915) );
  AN2 U2401 ( .A(n291), .B(n215), .Z(n1914) );
  AN2 U2402 ( .A(pos_disp_tx), .B(n81), .Z(n1913) );
  AN2 U2403 ( .A(n291), .B(n228), .Z(n1912) );
  AN2 U2404 ( .A(n291), .B(n277), .Z(n1911) );
  AN2 U2405 ( .A(n291), .B(n143), .Z(n1910) );
  AN2 U2406 ( .A(n291), .B(n191), .Z(n1909) );
  AN2 U2407 ( .A(n291), .B(n70), .Z(n1908) );
  AN2 U2408 ( .A(pos_disp_tx), .B(n241), .Z(n1907) );
  AN2 U2409 ( .A(pos_disp_tx), .B(n107), .Z(n1906) );
  AN2 U2410 ( .A(pos_disp_tx), .B(n58), .Z(n1905) );
  AN2 U2411 ( .A(n291), .B(n216), .Z(n1904) );
  AN2 U2412 ( .A(pos_disp_tx), .B(n82), .Z(n1903) );
  AN2 U2413 ( .A(n291), .B(n192), .Z(n1902) );
  AN2 U2414 ( .A(n291), .B(n71), .Z(n1901) );
  AN2 U2415 ( .A(n291), .B(n217), .Z(n1900) );
  AN2 U2416 ( .A(pos_disp_tx), .B(n83), .Z(n1899) );
  AN2 U2417 ( .A(n291), .B(n230), .Z(n1898) );
  AN2 U2418 ( .A(n291), .B(n279), .Z(n1897) );
  AN2 U2419 ( .A(n291), .B(n145), .Z(n1896) );
  AN2 U2420 ( .A(n291), .B(N239), .Z(n1895) );
  OR2 U2421 ( .A(n1893), .B(n1894), .Z(N835) );
  OR2 U2422 ( .A(n1891), .B(n1892), .Z(n1894) );
  OR2 U2423 ( .A(n1889), .B(n1890), .Z(n1893) );
  OR2 U2424 ( .A(n1887), .B(n1888), .Z(n1892) );
  OR2 U2425 ( .A(n1885), .B(n1886), .Z(n1891) );
  OR2 U2426 ( .A(n1883), .B(n1884), .Z(n1890) );
  OR2 U2427 ( .A(n1881), .B(n1882), .Z(n1889) );
  OR2 U2428 ( .A(n1880), .B(n1865), .Z(n1888) );
  OR2 U2429 ( .A(n1878), .B(n1879), .Z(n1887) );
  OR2 U2430 ( .A(n1876), .B(n1877), .Z(n1886) );
  OR2 U2431 ( .A(n1874), .B(n1875), .Z(n1885) );
  OR2 U2432 ( .A(n1872), .B(n1873), .Z(n1884) );
  OR2 U2433 ( .A(n1870), .B(n1871), .Z(n1883) );
  OR2 U2434 ( .A(n1868), .B(n1869), .Z(n1882) );
  OR2 U2435 ( .A(n1866), .B(n1867), .Z(n1881) );
  OR2 U2436 ( .A(n1863), .B(n1864), .Z(n1880) );
  OR2 U2437 ( .A(n1861), .B(n1862), .Z(n1879) );
  OR2 U2438 ( .A(n1859), .B(n1860), .Z(n1878) );
  OR2 U2439 ( .A(n1857), .B(n1858), .Z(n1877) );
  OR2 U2440 ( .A(n1855), .B(n1856), .Z(n1876) );
  OR2 U2441 ( .A(n1853), .B(n1854), .Z(n1875) );
  OR2 U2442 ( .A(n1851), .B(n1852), .Z(n1874) );
  OR2 U2443 ( .A(n1849), .B(n1850), .Z(n1873) );
  OR2 U2444 ( .A(n1847), .B(n1848), .Z(n1872) );
  OR2 U2445 ( .A(n1845), .B(n1846), .Z(n1871) );
  OR2 U2446 ( .A(n1843), .B(n1844), .Z(n1870) );
  OR2 U2447 ( .A(n1841), .B(n1842), .Z(n1869) );
  OR2 U2448 ( .A(n1839), .B(n1840), .Z(n1868) );
  OR2 U2449 ( .A(n1837), .B(n1838), .Z(n1867) );
  OR2 U2450 ( .A(n1835), .B(n1836), .Z(n1866) );
  OR2 U2451 ( .A(n1833), .B(n1834), .Z(n1865) );
  OR2 U2452 ( .A(n1831), .B(n1832), .Z(n1864) );
  OR2 U2453 ( .A(n1829), .B(n1830), .Z(n1863) );
  OR2 U2454 ( .A(n1827), .B(n1828), .Z(n1862) );
  OR2 U2455 ( .A(n1825), .B(n1826), .Z(n1861) );
  OR2 U2456 ( .A(n1823), .B(n1824), .Z(n1860) );
  OR2 U2457 ( .A(n1821), .B(n1822), .Z(n1859) );
  OR2 U2458 ( .A(n1819), .B(n1820), .Z(n1858) );
  OR2 U2459 ( .A(n1817), .B(n1818), .Z(n1857) );
  OR2 U2460 ( .A(n1815), .B(n1816), .Z(n1856) );
  OR2 U2461 ( .A(n1813), .B(n1814), .Z(n1855) );
  OR2 U2462 ( .A(n1811), .B(n1812), .Z(n1854) );
  OR2 U2463 ( .A(n1809), .B(n1810), .Z(n1853) );
  OR2 U2464 ( .A(n1807), .B(n1808), .Z(n1852) );
  OR2 U2465 ( .A(n1805), .B(n1806), .Z(n1851) );
  OR2 U2466 ( .A(n1803), .B(n1804), .Z(n1850) );
  OR2 U2467 ( .A(n1801), .B(n1802), .Z(n1849) );
  OR2 U2468 ( .A(n1799), .B(n1800), .Z(n1848) );
  OR2 U2469 ( .A(n1797), .B(n1798), .Z(n1847) );
  OR2 U2470 ( .A(n1795), .B(n1796), .Z(n1846) );
  OR2 U2471 ( .A(n1793), .B(n1794), .Z(n1845) );
  OR2 U2472 ( .A(n1791), .B(n1792), .Z(n1844) );
  OR2 U2473 ( .A(N955), .B(n1790), .Z(n1843) );
  OR2 U2474 ( .A(n1788), .B(n1789), .Z(n1842) );
  OR2 U2475 ( .A(n1786), .B(n1787), .Z(n1841) );
  OR2 U2476 ( .A(n1784), .B(n1785), .Z(n1840) );
  OR2 U2477 ( .A(n1782), .B(n1783), .Z(n1839) );
  OR2 U2478 ( .A(n1780), .B(n1781), .Z(n1838) );
  OR2 U2479 ( .A(n1778), .B(n1779), .Z(n1837) );
  OR2 U2480 ( .A(n1776), .B(n1777), .Z(n1836) );
  OR2 U2481 ( .A(n1774), .B(n1775), .Z(n1835) );
  OR2 U2482 ( .A(n1772), .B(n1773), .Z(n1834) );
  OR2 U2483 ( .A(n1770), .B(n1771), .Z(n1833) );
  OR2 U2484 ( .A(n1768), .B(n1769), .Z(n1832) );
  OR2 U2485 ( .A(n1766), .B(n1767), .Z(n1831) );
  OR2 U2486 ( .A(n1764), .B(n1765), .Z(n1830) );
  OR2 U2487 ( .A(n1762), .B(n1763), .Z(n1829) );
  OR2 U2488 ( .A(n1760), .B(n1761), .Z(n1828) );
  OR2 U2489 ( .A(n1758), .B(n1759), .Z(n1827) );
  OR2 U2490 ( .A(n1756), .B(n1757), .Z(n1826) );
  OR2 U2491 ( .A(n1754), .B(n1755), .Z(n1825) );
  OR2 U2492 ( .A(n1752), .B(n1753), .Z(n1824) );
  OR2 U2493 ( .A(n1750), .B(n1751), .Z(n1823) );
  OR2 U2494 ( .A(n1748), .B(n1749), .Z(n1822) );
  OR2 U2495 ( .A(n1746), .B(n1747), .Z(n1821) );
  OR2 U2496 ( .A(n1744), .B(n1745), .Z(n1820) );
  OR2 U2497 ( .A(n1742), .B(n1743), .Z(n1819) );
  OR2 U2498 ( .A(n1740), .B(n1741), .Z(n1818) );
  OR2 U2499 ( .A(n1738), .B(n1739), .Z(n1817) );
  OR2 U2500 ( .A(n1736), .B(n1737), .Z(n1816) );
  OR2 U2501 ( .A(n1734), .B(n1735), .Z(n1815) );
  OR2 U2502 ( .A(n1732), .B(n1733), .Z(n1814) );
  OR2 U2503 ( .A(n1730), .B(n1731), .Z(n1813) );
  OR2 U2504 ( .A(n1728), .B(n1729), .Z(n1812) );
  OR2 U2505 ( .A(n1726), .B(n1727), .Z(n1811) );
  OR2 U2506 ( .A(n1724), .B(n1725), .Z(n1810) );
  OR2 U2507 ( .A(n1722), .B(n1723), .Z(n1809) );
  OR2 U2508 ( .A(n1720), .B(n1721), .Z(n1808) );
  OR2 U2509 ( .A(n1718), .B(n1719), .Z(n1807) );
  OR2 U2510 ( .A(n1716), .B(n1717), .Z(n1806) );
  OR2 U2511 ( .A(n1714), .B(n1715), .Z(n1805) );
  OR2 U2512 ( .A(n1712), .B(n1713), .Z(n1804) );
  OR2 U2513 ( .A(n1710), .B(n1711), .Z(n1803) );
  OR2 U2514 ( .A(n1708), .B(n1709), .Z(n1802) );
  OR2 U2515 ( .A(n1706), .B(n1707), .Z(n1801) );
  OR2 U2516 ( .A(n1704), .B(n1705), .Z(n1800) );
  OR2 U2517 ( .A(n1702), .B(n1703), .Z(n1799) );
  OR2 U2518 ( .A(n1700), .B(n1701), .Z(n1798) );
  OR2 U2519 ( .A(n1698), .B(n1699), .Z(n1797) );
  OR2 U2520 ( .A(n1696), .B(n1697), .Z(n1796) );
  OR2 U2521 ( .A(n1694), .B(n1695), .Z(n1795) );
  OR2 U2522 ( .A(n1692), .B(n1693), .Z(n1794) );
  OR2 U2523 ( .A(n1690), .B(n1691), .Z(n1793) );
  OR2 U2524 ( .A(n1688), .B(n1689), .Z(n1792) );
  OR2 U2525 ( .A(n1686), .B(n1687), .Z(n1791) );
  OR2 U2526 ( .A(n1684), .B(n1685), .Z(n1790) );
  OR2 U2527 ( .A(n1682), .B(n1683), .Z(n1789) );
  OR2 U2528 ( .A(n1680), .B(n1681), .Z(n1788) );
  OR2 U2529 ( .A(n1678), .B(n1679), .Z(n1787) );
  OR2 U2530 ( .A(n1676), .B(n1677), .Z(n1786) );
  OR2 U2531 ( .A(n1674), .B(n1675), .Z(n1785) );
  OR2 U2532 ( .A(n1672), .B(n1673), .Z(n1784) );
  OR2 U2533 ( .A(n1670), .B(n1671), .Z(n1783) );
  OR2 U2534 ( .A(n1668), .B(n1669), .Z(n1782) );
  OR2 U2535 ( .A(n1666), .B(n1667), .Z(n1781) );
  OR2 U2536 ( .A(n1664), .B(n1665), .Z(n1780) );
  OR2 U2537 ( .A(n1662), .B(n1663), .Z(n1779) );
  OR2 U2538 ( .A(n1660), .B(n1661), .Z(n1778) );
  OR2 U2539 ( .A(n1658), .B(n1659), .Z(n1777) );
  OR2 U2540 ( .A(n1656), .B(n1657), .Z(n1776) );
  OR2 U2541 ( .A(n1654), .B(n1655), .Z(n1775) );
  OR2 U2542 ( .A(n1652), .B(n1653), .Z(n1774) );
  AN2 U2543 ( .A(pos_disp_tx), .B(N8311), .Z(n1773) );
  AN2 U2544 ( .A(pos_disp_tx), .B(n153), .Z(n1772) );
  AN2 U2545 ( .A(pos_disp_tx), .B(n33), .Z(n1771) );
  AN2 U2546 ( .A(n291), .B(n168), .Z(n1770) );
  AN2 U2547 ( .A(pos_disp_tx), .B(n19), .Z(n1769) );
  AN2 U2548 ( .A(n291), .B(n157), .Z(n1768) );
  AN2 U2549 ( .A(n291), .B(n37), .Z(n1767) );
  AN2 U2550 ( .A(pos_disp_tx), .B(n172), .Z(n1766) );
  AN2 U2551 ( .A(pos_disp_tx), .B(n26), .Z(n1765) );
  AN2 U2552 ( .A(n291), .B(n161), .Z(n1764) );
  AN2 U2553 ( .A(n291), .B(n40), .Z(n1763) );
  AN2 U2554 ( .A(n291), .B(n30), .Z(n1762) );
  AN2 U2555 ( .A(pos_disp_tx), .B(n178), .Z(n1761) );
  AN2 U2556 ( .A(pos_disp_tx), .B(n23), .Z(n1760) );
  AN2 U2557 ( .A(n291), .B(n169), .Z(n1759) );
  AN2 U2558 ( .A(n291), .B(n158), .Z(n1758) );
  AN2 U2559 ( .A(n291), .B(n38), .Z(n1757) );
  AN2 U2560 ( .A(pos_disp_tx), .B(n173), .Z(n1756) );
  AN2 U2561 ( .A(n291), .B(n27), .Z(n1755) );
  AN2 U2562 ( .A(n291), .B(n162), .Z(n1754) );
  AN2 U2563 ( .A(n291), .B(n41), .Z(n1753) );
  AN2 U2564 ( .A(pos_disp_tx), .B(n176), .Z(n1752) );
  AN2 U2565 ( .A(n291), .B(n31), .Z(n1751) );
  AN2 U2566 ( .A(pos_disp_tx), .B(n166), .Z(n1750) );
  AN2 U2567 ( .A(pos_disp_tx), .B(n44), .Z(n1749) );
  AN2 U2568 ( .A(pos_disp_tx), .B(n179), .Z(n1748) );
  AN2 U2569 ( .A(pos_disp_tx), .B(n62), .Z(n1747) );
  AN2 U2570 ( .A(pos_disp_tx), .B(n233), .Z(n1746) );
  AN2 U2571 ( .A(pos_disp_tx), .B(n99), .Z(n1745) );
  AN2 U2572 ( .A(n291), .B(n195), .Z(n1744) );
  AN2 U2573 ( .A(pos_disp_tx), .B(n50), .Z(n1743) );
  AN2 U2574 ( .A(n291), .B(n245), .Z(n1742) );
  AN2 U2575 ( .A(n291), .B(n111), .Z(n1741) );
  AN2 U2576 ( .A(pos_disp_tx), .B(n208), .Z(n1740) );
  AN2 U2577 ( .A(pos_disp_tx), .B(n74), .Z(n1739) );
  AN2 U2578 ( .A(n291), .B(n257), .Z(n1738) );
  AN2 U2579 ( .A(n291), .B(n123), .Z(n1737) );
  AN2 U2580 ( .A(n291), .B(n221), .Z(n1736) );
  AN2 U2581 ( .A(n291), .B(n87), .Z(n1735) );
  AN2 U2582 ( .A(n291), .B(n270), .Z(n1734) );
  AN2 U2583 ( .A(n291), .B(n136), .Z(n1733) );
  AN2 U2584 ( .A(pos_disp_tx), .B(n184), .Z(n1732) );
  AN2 U2585 ( .A(pos_disp_tx), .B(n63), .Z(n1731) );
  AN2 U2586 ( .A(n291), .B(n234), .Z(n1730) );
  AN2 U2587 ( .A(n291), .B(n100), .Z(n1729) );
  AN2 U2588 ( .A(n291), .B(n196), .Z(n1728) );
  AN2 U2589 ( .A(n291), .B(n51), .Z(n1727) );
  AN2 U2590 ( .A(n291), .B(n246), .Z(n1726) );
  AN2 U2591 ( .A(n291), .B(n112), .Z(n1725) );
  AN2 U2592 ( .A(pos_disp_tx), .B(n209), .Z(n1724) );
  AN2 U2593 ( .A(n291), .B(n75), .Z(n1723) );
  AN2 U2594 ( .A(n291), .B(n258), .Z(n1722) );
  AN2 U2595 ( .A(n291), .B(n124), .Z(n1721) );
  AN2 U2596 ( .A(pos_disp_tx), .B(n222), .Z(n1720) );
  AN2 U2597 ( .A(n291), .B(n88), .Z(n1719) );
  AN2 U2598 ( .A(pos_disp_tx), .B(n271), .Z(n1718) );
  AN2 U2599 ( .A(pos_disp_tx), .B(n137), .Z(n1717) );
  AN2 U2600 ( .A(pos_disp_tx), .B(n185), .Z(n1716) );
  AN2 U2601 ( .A(pos_disp_tx), .B(n64), .Z(n1715) );
  AN2 U2602 ( .A(pos_disp_tx), .B(n235), .Z(n1714) );
  AN2 U2603 ( .A(pos_disp_tx), .B(n101), .Z(n1713) );
  AN2 U2604 ( .A(n291), .B(n197), .Z(n1712) );
  AN2 U2605 ( .A(pos_disp_tx), .B(n52), .Z(n1711) );
  AN2 U2606 ( .A(n291), .B(n247), .Z(n1710) );
  AN2 U2607 ( .A(n291), .B(n113), .Z(n1709) );
  AN2 U2608 ( .A(pos_disp_tx), .B(n210), .Z(n1708) );
  AN2 U2609 ( .A(pos_disp_tx), .B(n76), .Z(n1707) );
  AN2 U2610 ( .A(n291), .B(n259), .Z(n1706) );
  AN2 U2611 ( .A(n291), .B(n125), .Z(n1705) );
  AN2 U2612 ( .A(n291), .B(n223), .Z(n1704) );
  AN2 U2613 ( .A(n291), .B(n89), .Z(n1703) );
  AN2 U2614 ( .A(n291), .B(n272), .Z(n1702) );
  AN2 U2615 ( .A(n291), .B(n138), .Z(n1701) );
  AN2 U2616 ( .A(pos_disp_tx), .B(n186), .Z(n1700) );
  AN2 U2617 ( .A(pos_disp_tx), .B(n65), .Z(n1699) );
  AN2 U2618 ( .A(n291), .B(n236), .Z(n1698) );
  AN2 U2619 ( .A(n291), .B(n102), .Z(n1697) );
  AN2 U2620 ( .A(n291), .B(n198), .Z(n1696) );
  AN2 U2621 ( .A(n291), .B(n53), .Z(n1695) );
  AN2 U2622 ( .A(n291), .B(n248), .Z(n1694) );
  AN2 U2623 ( .A(n291), .B(n114), .Z(n1693) );
  AN2 U2624 ( .A(pos_disp_tx), .B(n211), .Z(n1692) );
  AN2 U2625 ( .A(n291), .B(n77), .Z(n1691) );
  AN2 U2626 ( .A(n291), .B(n260), .Z(n1690) );
  AN2 U2627 ( .A(n291), .B(n126), .Z(n1689) );
  AN2 U2628 ( .A(pos_disp_tx), .B(n224), .Z(n1688) );
  AN2 U2629 ( .A(n291), .B(n90), .Z(n1687) );
  AN2 U2630 ( .A(pos_disp_tx), .B(n273), .Z(n1686) );
  AN2 U2631 ( .A(pos_disp_tx), .B(n139), .Z(n1685) );
  AN2 U2632 ( .A(pos_disp_tx), .B(n187), .Z(n1684) );
  AN2 U2633 ( .A(pos_disp_tx), .B(n70), .Z(n1683) );
  AN2 U2634 ( .A(pos_disp_tx), .B(n241), .Z(n1682) );
  AN2 U2635 ( .A(pos_disp_tx), .B(n107), .Z(n1681) );
  AN2 U2636 ( .A(n291), .B(n203), .Z(n1680) );
  AN2 U2637 ( .A(pos_disp_tx), .B(n58), .Z(n1679) );
  AN2 U2638 ( .A(n291), .B(n253), .Z(n1678) );
  AN2 U2639 ( .A(n291), .B(n119), .Z(n1677) );
  AN2 U2640 ( .A(pos_disp_tx), .B(n216), .Z(n1676) );
  AN2 U2641 ( .A(pos_disp_tx), .B(n82), .Z(n1675) );
  AN2 U2642 ( .A(n291), .B(n265), .Z(n1674) );
  AN2 U2643 ( .A(n291), .B(n131), .Z(n1673) );
  AN2 U2644 ( .A(n291), .B(n229), .Z(n1672) );
  AN2 U2645 ( .A(n291), .B(n95), .Z(n1671) );
  AN2 U2646 ( .A(n291), .B(n278), .Z(n1670) );
  AN2 U2647 ( .A(n291), .B(n144), .Z(n1669) );
  AN2 U2648 ( .A(pos_disp_tx), .B(n192), .Z(n1668) );
  AN2 U2649 ( .A(pos_disp_tx), .B(n71), .Z(n1667) );
  AN2 U2650 ( .A(n291), .B(n242), .Z(n1666) );
  AN2 U2651 ( .A(n291), .B(n108), .Z(n1665) );
  AN2 U2652 ( .A(n291), .B(n204), .Z(n1664) );
  AN2 U2653 ( .A(n291), .B(n59), .Z(n1663) );
  AN2 U2654 ( .A(n291), .B(n254), .Z(n1662) );
  AN2 U2655 ( .A(n291), .B(n120), .Z(n1661) );
  AN2 U2656 ( .A(pos_disp_tx), .B(n217), .Z(n1660) );
  AN2 U2657 ( .A(n291), .B(n83), .Z(n1659) );
  AN2 U2658 ( .A(n291), .B(n266), .Z(n1658) );
  AN2 U2659 ( .A(n291), .B(n132), .Z(n1657) );
  AN2 U2660 ( .A(pos_disp_tx), .B(n230), .Z(n1656) );
  AN2 U2661 ( .A(n291), .B(n96), .Z(n1655) );
  AN2 U2662 ( .A(pos_disp_tx), .B(n279), .Z(n1654) );
  AN2 U2663 ( .A(pos_disp_tx), .B(n145), .Z(n1653) );
  AN2 U2664 ( .A(pos_disp_tx), .B(N239), .Z(n1652) );
  OR2 U2665 ( .A(n1651), .B(n1588), .Z(N834) );
  OR2 U2666 ( .A(n1649), .B(n1650), .Z(n1651) );
  OR2 U2667 ( .A(n1647), .B(n1648), .Z(n1650) );
  OR2 U2668 ( .A(n1645), .B(n1646), .Z(n1649) );
  OR2 U2669 ( .A(n1643), .B(n1644), .Z(n1648) );
  OR2 U2670 ( .A(n1641), .B(n1642), .Z(n1647) );
  OR2 U2671 ( .A(n1639), .B(n1640), .Z(n1646) );
  OR2 U2672 ( .A(n1637), .B(n1638), .Z(n1645) );
  OR2 U2673 ( .A(n1635), .B(n1636), .Z(n1644) );
  OR2 U2674 ( .A(n1633), .B(n1634), .Z(n1643) );
  OR2 U2675 ( .A(n1631), .B(n1632), .Z(n1642) );
  OR2 U2676 ( .A(n1629), .B(n1630), .Z(n1641) );
  OR2 U2677 ( .A(n1627), .B(n1628), .Z(n1640) );
  OR2 U2678 ( .A(n1625), .B(n1626), .Z(n1639) );
  OR2 U2679 ( .A(n1623), .B(n1624), .Z(n1638) );
  OR2 U2680 ( .A(n1621), .B(n1622), .Z(n1637) );
  OR2 U2681 ( .A(n1619), .B(n1620), .Z(n1636) );
  OR2 U2682 ( .A(n1617), .B(n1618), .Z(n1635) );
  OR2 U2683 ( .A(n1615), .B(n1616), .Z(n1634) );
  OR2 U2684 ( .A(n1613), .B(n1614), .Z(n1633) );
  OR2 U2685 ( .A(n1611), .B(n1612), .Z(n1632) );
  OR2 U2686 ( .A(n1609), .B(n1610), .Z(n1631) );
  OR2 U2687 ( .A(n1607), .B(n1608), .Z(n1630) );
  OR2 U2688 ( .A(n1605), .B(n1606), .Z(n1629) );
  OR2 U2689 ( .A(n1603), .B(n1604), .Z(n1628) );
  OR2 U2690 ( .A(n1601), .B(n1602), .Z(n1627) );
  OR2 U2691 ( .A(n1599), .B(n1600), .Z(n1626) );
  OR2 U2692 ( .A(n1597), .B(n1598), .Z(n1625) );
  OR2 U2693 ( .A(n1595), .B(n1596), .Z(n1624) );
  OR2 U2694 ( .A(n1593), .B(n1594), .Z(n1623) );
  OR2 U2695 ( .A(n1591), .B(n1592), .Z(n1622) );
  OR2 U2696 ( .A(n1589), .B(n1590), .Z(n1621) );
  OR2 U2697 ( .A(n1586), .B(n1587), .Z(n1620) );
  OR2 U2698 ( .A(n1584), .B(n1585), .Z(n1619) );
  OR2 U2699 ( .A(n1582), .B(n1583), .Z(n1618) );
  OR2 U2700 ( .A(n1580), .B(n1581), .Z(n1617) );
  OR2 U2701 ( .A(n1578), .B(n1579), .Z(n1616) );
  OR2 U2702 ( .A(n1576), .B(n1577), .Z(n1615) );
  OR2 U2703 ( .A(n1574), .B(n1575), .Z(n1614) );
  OR2 U2704 ( .A(n1572), .B(n1573), .Z(n1613) );
  OR2 U2705 ( .A(n1570), .B(n1571), .Z(n1612) );
  OR2 U2706 ( .A(n1568), .B(n1569), .Z(n1611) );
  OR2 U2707 ( .A(n1566), .B(n1567), .Z(n1610) );
  OR2 U2708 ( .A(n1564), .B(n1565), .Z(n1609) );
  OR2 U2709 ( .A(n1562), .B(n1563), .Z(n1608) );
  OR2 U2710 ( .A(n1560), .B(n1561), .Z(n1607) );
  OR2 U2711 ( .A(n1558), .B(n1559), .Z(n1606) );
  OR2 U2712 ( .A(n1556), .B(n1557), .Z(n1605) );
  OR2 U2713 ( .A(n1554), .B(n1555), .Z(n1604) );
  OR2 U2714 ( .A(n1552), .B(n1553), .Z(n1603) );
  OR2 U2715 ( .A(n1550), .B(n1551), .Z(n1602) );
  OR2 U2716 ( .A(n1548), .B(n1549), .Z(n1601) );
  OR2 U2717 ( .A(n1546), .B(n1547), .Z(n1600) );
  OR2 U2718 ( .A(n1544), .B(n1545), .Z(n1599) );
  OR2 U2719 ( .A(n1542), .B(n1543), .Z(n1598) );
  OR2 U2720 ( .A(N952), .B(n1541), .Z(n1597) );
  OR2 U2721 ( .A(n1539), .B(n1540), .Z(n1596) );
  OR2 U2722 ( .A(n1537), .B(n1538), .Z(n1595) );
  OR2 U2723 ( .A(n1535), .B(n1536), .Z(n1594) );
  OR2 U2724 ( .A(n1533), .B(n1534), .Z(n1593) );
  OR2 U2725 ( .A(n1531), .B(n1532), .Z(n1592) );
  OR2 U2726 ( .A(n1529), .B(n1530), .Z(n1591) );
  OR2 U2727 ( .A(n1527), .B(n1528), .Z(n1590) );
  OR2 U2728 ( .A(n1525), .B(n1526), .Z(n1589) );
  OR2 U2729 ( .A(n1523), .B(n1524), .Z(n1588) );
  OR2 U2730 ( .A(n1521), .B(n1522), .Z(n1587) );
  OR2 U2731 ( .A(n1519), .B(n1520), .Z(n1586) );
  OR2 U2732 ( .A(n1517), .B(n1518), .Z(n1585) );
  OR2 U2733 ( .A(n1515), .B(n1516), .Z(n1584) );
  OR2 U2734 ( .A(n1513), .B(n1514), .Z(n1583) );
  OR2 U2735 ( .A(n1511), .B(n1512), .Z(n1582) );
  OR2 U2736 ( .A(n1509), .B(n1510), .Z(n1581) );
  OR2 U2737 ( .A(n1507), .B(n1508), .Z(n1580) );
  OR2 U2738 ( .A(n1505), .B(n1506), .Z(n1579) );
  OR2 U2739 ( .A(n1503), .B(n1504), .Z(n1578) );
  OR2 U2740 ( .A(n1501), .B(n1502), .Z(n1577) );
  OR2 U2741 ( .A(n1499), .B(n1500), .Z(n1576) );
  OR2 U2742 ( .A(n1497), .B(n1498), .Z(n1575) );
  OR2 U2743 ( .A(n1495), .B(n1496), .Z(n1574) );
  OR2 U2744 ( .A(n1493), .B(n1494), .Z(n1573) );
  OR2 U2745 ( .A(n1491), .B(n1492), .Z(n1572) );
  OR2 U2746 ( .A(n1489), .B(n1490), .Z(n1571) );
  OR2 U2747 ( .A(n1487), .B(n1488), .Z(n1570) );
  OR2 U2748 ( .A(n1485), .B(n1486), .Z(n1569) );
  OR2 U2749 ( .A(n1483), .B(n1484), .Z(n1568) );
  OR2 U2750 ( .A(n1481), .B(n1482), .Z(n1567) );
  OR2 U2751 ( .A(n1479), .B(n1480), .Z(n1566) );
  OR2 U2752 ( .A(n1477), .B(n1478), .Z(n1565) );
  OR2 U2753 ( .A(n1475), .B(n1476), .Z(n1564) );
  OR2 U2754 ( .A(n1473), .B(n1474), .Z(n1563) );
  OR2 U2755 ( .A(n1471), .B(n1472), .Z(n1562) );
  OR2 U2756 ( .A(n1469), .B(n1470), .Z(n1561) );
  OR2 U2757 ( .A(n1467), .B(n1468), .Z(n1560) );
  OR2 U2758 ( .A(n1465), .B(n1466), .Z(n1559) );
  OR2 U2759 ( .A(n1463), .B(n1464), .Z(n1558) );
  OR2 U2760 ( .A(n1461), .B(n1462), .Z(n1557) );
  OR2 U2761 ( .A(n1459), .B(n1460), .Z(n1556) );
  OR2 U2762 ( .A(n1457), .B(n1458), .Z(n1555) );
  OR2 U2763 ( .A(n1455), .B(n1456), .Z(n1554) );
  OR2 U2764 ( .A(n1453), .B(n1454), .Z(n1553) );
  OR2 U2765 ( .A(n1451), .B(n1452), .Z(n1552) );
  OR2 U2766 ( .A(n1449), .B(n1450), .Z(n1551) );
  OR2 U2767 ( .A(n1447), .B(n1448), .Z(n1550) );
  OR2 U2768 ( .A(n1445), .B(n1446), .Z(n1549) );
  OR2 U2769 ( .A(n1443), .B(n1444), .Z(n1548) );
  OR2 U2770 ( .A(n1441), .B(n1442), .Z(n1547) );
  OR2 U2771 ( .A(n1439), .B(n1440), .Z(n1546) );
  OR2 U2772 ( .A(n1437), .B(n1438), .Z(n1545) );
  OR2 U2773 ( .A(n1435), .B(n1436), .Z(n1544) );
  OR2 U2774 ( .A(n1433), .B(n1434), .Z(n1543) );
  OR2 U2775 ( .A(n1431), .B(n1432), .Z(n1542) );
  OR2 U2776 ( .A(n1429), .B(n1430), .Z(n1541) );
  OR2 U2777 ( .A(n1427), .B(n1428), .Z(n1540) );
  OR2 U2778 ( .A(n1425), .B(n1426), .Z(n1539) );
  OR2 U2779 ( .A(n1423), .B(n1424), .Z(n1538) );
  OR2 U2780 ( .A(n1421), .B(n1422), .Z(n1537) );
  OR2 U2781 ( .A(n1419), .B(n1420), .Z(n1536) );
  OR2 U2782 ( .A(n1417), .B(n1418), .Z(n1535) );
  OR2 U2783 ( .A(n1415), .B(n1416), .Z(n1534) );
  OR2 U2784 ( .A(n1413), .B(n1414), .Z(n1533) );
  OR2 U2785 ( .A(n1411), .B(n1412), .Z(n1532) );
  OR2 U2786 ( .A(n1409), .B(n1410), .Z(n1531) );
  OR2 U2787 ( .A(n1407), .B(n1408), .Z(n1530) );
  OR2 U2788 ( .A(n1405), .B(n1406), .Z(n1529) );
  OR2 U2789 ( .A(n1403), .B(n1404), .Z(n1528) );
  OR2 U2790 ( .A(n1401), .B(n1402), .Z(n1527) );
  OR2 U2791 ( .A(n1399), .B(n1400), .Z(n1526) );
  OR2 U2792 ( .A(n1397), .B(n1398), .Z(n1525) );
  AN2 U2793 ( .A(pos_disp_tx), .B(N8311), .Z(n1524) );
  AN2 U2794 ( .A(pos_disp_tx), .B(n153), .Z(n1523) );
  AN2 U2795 ( .A(pos_disp_tx), .B(n33), .Z(n1522) );
  AN2 U2796 ( .A(n291), .B(n168), .Z(n1521) );
  AN2 U2797 ( .A(pos_disp_tx), .B(n19), .Z(n1520) );
  AN2 U2798 ( .A(n291), .B(n157), .Z(n1519) );
  AN2 U2799 ( .A(n291), .B(n37), .Z(n1518) );
  AN2 U2800 ( .A(pos_disp_tx), .B(n172), .Z(n1517) );
  AN2 U2801 ( .A(pos_disp_tx), .B(n26), .Z(n1516) );
  AN2 U2802 ( .A(n291), .B(n161), .Z(n1515) );
  AN2 U2803 ( .A(n291), .B(n40), .Z(n1514) );
  AN2 U2804 ( .A(n291), .B(n175), .Z(n1513) );
  AN2 U2805 ( .A(n291), .B(n30), .Z(n1512) );
  AN2 U2806 ( .A(n291), .B(n165), .Z(n1511) );
  AN2 U2807 ( .A(n291), .B(n43), .Z(n1510) );
  AN2 U2808 ( .A(pos_disp_tx), .B(n178), .Z(n1509) );
  AN2 U2809 ( .A(pos_disp_tx), .B(n23), .Z(n1508) );
  AN2 U2810 ( .A(n291), .B(n154), .Z(n1507) );
  AN2 U2811 ( .A(n291), .B(n34), .Z(n1506) );
  AN2 U2812 ( .A(n291), .B(n169), .Z(n1505) );
  AN2 U2813 ( .A(n291), .B(n20), .Z(n1504) );
  AN2 U2814 ( .A(n291), .B(n158), .Z(n1503) );
  AN2 U2815 ( .A(n291), .B(n38), .Z(n1502) );
  AN2 U2816 ( .A(pos_disp_tx), .B(n173), .Z(n1501) );
  AN2 U2817 ( .A(n291), .B(n27), .Z(n1500) );
  AN2 U2818 ( .A(n291), .B(n162), .Z(n1499) );
  AN2 U2819 ( .A(n291), .B(n41), .Z(n1498) );
  AN2 U2820 ( .A(pos_disp_tx), .B(n176), .Z(n1497) );
  AN2 U2821 ( .A(n291), .B(n31), .Z(n1496) );
  AN2 U2822 ( .A(pos_disp_tx), .B(n166), .Z(n1495) );
  AN2 U2823 ( .A(pos_disp_tx), .B(n44), .Z(n1494) );
  AN2 U2824 ( .A(pos_disp_tx), .B(n179), .Z(n1493) );
  AN2 U2825 ( .A(pos_disp_tx), .B(n62), .Z(n1492) );
  AN2 U2826 ( .A(pos_disp_tx), .B(n233), .Z(n1491) );
  AN2 U2827 ( .A(pos_disp_tx), .B(n99), .Z(n1490) );
  AN2 U2828 ( .A(n291), .B(n195), .Z(n1489) );
  AN2 U2829 ( .A(pos_disp_tx), .B(n50), .Z(n1488) );
  AN2 U2830 ( .A(n291), .B(n245), .Z(n1487) );
  AN2 U2831 ( .A(n291), .B(n111), .Z(n1486) );
  AN2 U2832 ( .A(pos_disp_tx), .B(n208), .Z(n1485) );
  AN2 U2833 ( .A(pos_disp_tx), .B(n74), .Z(n1484) );
  AN2 U2834 ( .A(n291), .B(n257), .Z(n1483) );
  AN2 U2835 ( .A(n291), .B(n123), .Z(n1482) );
  AN2 U2836 ( .A(n291), .B(n221), .Z(n1481) );
  AN2 U2837 ( .A(n291), .B(n87), .Z(n1480) );
  AN2 U2838 ( .A(n291), .B(n270), .Z(n1479) );
  AN2 U2839 ( .A(n291), .B(n136), .Z(n1478) );
  AN2 U2840 ( .A(pos_disp_tx), .B(n184), .Z(n1477) );
  AN2 U2841 ( .A(pos_disp_tx), .B(n63), .Z(n1476) );
  AN2 U2842 ( .A(n291), .B(n234), .Z(n1475) );
  AN2 U2843 ( .A(n291), .B(n100), .Z(n1474) );
  AN2 U2844 ( .A(n291), .B(n196), .Z(n1473) );
  AN2 U2845 ( .A(n291), .B(n51), .Z(n1472) );
  AN2 U2846 ( .A(n291), .B(n246), .Z(n1471) );
  AN2 U2847 ( .A(n291), .B(n112), .Z(n1470) );
  AN2 U2848 ( .A(pos_disp_tx), .B(n209), .Z(n1469) );
  AN2 U2849 ( .A(n291), .B(n75), .Z(n1468) );
  AN2 U2850 ( .A(n291), .B(n258), .Z(n1467) );
  AN2 U2851 ( .A(n291), .B(n124), .Z(n1466) );
  AN2 U2852 ( .A(pos_disp_tx), .B(n222), .Z(n1465) );
  AN2 U2853 ( .A(n291), .B(n88), .Z(n1464) );
  AN2 U2854 ( .A(pos_disp_tx), .B(n271), .Z(n1463) );
  AN2 U2855 ( .A(pos_disp_tx), .B(n137), .Z(n1462) );
  AN2 U2856 ( .A(pos_disp_tx), .B(n185), .Z(n1461) );
  AN2 U2857 ( .A(pos_disp_tx), .B(n64), .Z(n1460) );
  AN2 U2858 ( .A(pos_disp_tx), .B(n235), .Z(n1459) );
  AN2 U2859 ( .A(pos_disp_tx), .B(n101), .Z(n1458) );
  AN2 U2860 ( .A(n291), .B(n197), .Z(n1457) );
  AN2 U2861 ( .A(pos_disp_tx), .B(n52), .Z(n1456) );
  AN2 U2862 ( .A(n291), .B(n247), .Z(n1455) );
  AN2 U2863 ( .A(n291), .B(n113), .Z(n1454) );
  AN2 U2864 ( .A(pos_disp_tx), .B(n210), .Z(n1453) );
  AN2 U2865 ( .A(pos_disp_tx), .B(n76), .Z(n1452) );
  AN2 U2866 ( .A(n291), .B(n259), .Z(n1451) );
  AN2 U2867 ( .A(n291), .B(n125), .Z(n1450) );
  AN2 U2868 ( .A(n291), .B(n223), .Z(n1449) );
  AN2 U2869 ( .A(n291), .B(n89), .Z(n1448) );
  AN2 U2870 ( .A(n291), .B(n272), .Z(n1447) );
  AN2 U2871 ( .A(n291), .B(n138), .Z(n1446) );
  AN2 U2872 ( .A(pos_disp_tx), .B(n186), .Z(n1445) );
  AN2 U2873 ( .A(pos_disp_tx), .B(n65), .Z(n1444) );
  AN2 U2874 ( .A(n291), .B(n236), .Z(n1443) );
  AN2 U2875 ( .A(n291), .B(n102), .Z(n1442) );
  AN2 U2876 ( .A(n291), .B(n198), .Z(n1441) );
  AN2 U2877 ( .A(n291), .B(n53), .Z(n1440) );
  AN2 U2878 ( .A(n291), .B(n248), .Z(n1439) );
  AN2 U2879 ( .A(n291), .B(n114), .Z(n1438) );
  AN2 U2880 ( .A(pos_disp_tx), .B(n211), .Z(n1437) );
  AN2 U2881 ( .A(n291), .B(n77), .Z(n1436) );
  AN2 U2882 ( .A(n291), .B(n260), .Z(n1435) );
  AN2 U2883 ( .A(n291), .B(n126), .Z(n1434) );
  AN2 U2884 ( .A(pos_disp_tx), .B(n224), .Z(n1433) );
  AN2 U2885 ( .A(n291), .B(n90), .Z(n1432) );
  AN2 U2886 ( .A(pos_disp_tx), .B(n273), .Z(n1431) );
  AN2 U2887 ( .A(pos_disp_tx), .B(n139), .Z(n1430) );
  AN2 U2888 ( .A(pos_disp_tx), .B(n187), .Z(n1429) );
  AN2 U2889 ( .A(n291), .B(n70), .Z(n1428) );
  AN2 U2890 ( .A(n291), .B(n241), .Z(n1427) );
  AN2 U2891 ( .A(n291), .B(n107), .Z(n1426) );
  AN2 U2892 ( .A(pos_disp_tx), .B(n203), .Z(n1425) );
  AN2 U2893 ( .A(n291), .B(n58), .Z(n1424) );
  AN2 U2894 ( .A(pos_disp_tx), .B(n253), .Z(n1423) );
  AN2 U2895 ( .A(pos_disp_tx), .B(n119), .Z(n1422) );
  AN2 U2896 ( .A(n291), .B(n216), .Z(n1421) );
  AN2 U2897 ( .A(n291), .B(n82), .Z(n1420) );
  AN2 U2898 ( .A(pos_disp_tx), .B(n265), .Z(n1419) );
  AN2 U2899 ( .A(pos_disp_tx), .B(n131), .Z(n1418) );
  AN2 U2900 ( .A(pos_disp_tx), .B(n229), .Z(n1417) );
  AN2 U2901 ( .A(pos_disp_tx), .B(n95), .Z(n1416) );
  AN2 U2902 ( .A(pos_disp_tx), .B(n278), .Z(n1415) );
  AN2 U2903 ( .A(pos_disp_tx), .B(n144), .Z(n1414) );
  AN2 U2904 ( .A(n291), .B(n192), .Z(n1413) );
  AN2 U2905 ( .A(n291), .B(n71), .Z(n1412) );
  AN2 U2906 ( .A(pos_disp_tx), .B(n242), .Z(n1411) );
  AN2 U2907 ( .A(pos_disp_tx), .B(n108), .Z(n1410) );
  AN2 U2908 ( .A(pos_disp_tx), .B(n204), .Z(n1409) );
  AN2 U2909 ( .A(pos_disp_tx), .B(n59), .Z(n1408) );
  AN2 U2910 ( .A(pos_disp_tx), .B(n254), .Z(n1407) );
  AN2 U2911 ( .A(pos_disp_tx), .B(n120), .Z(n1406) );
  AN2 U2912 ( .A(n291), .B(n217), .Z(n1405) );
  AN2 U2913 ( .A(pos_disp_tx), .B(n83), .Z(n1404) );
  AN2 U2914 ( .A(pos_disp_tx), .B(n266), .Z(n1403) );
  AN2 U2915 ( .A(pos_disp_tx), .B(n132), .Z(n1402) );
  AN2 U2916 ( .A(n291), .B(n230), .Z(n1401) );
  AN2 U2917 ( .A(pos_disp_tx), .B(n96), .Z(n1400) );
  AN2 U2918 ( .A(n291), .B(n279), .Z(n1399) );
  AN2 U2919 ( .A(n291), .B(n145), .Z(n1398) );
  AN2 U2920 ( .A(n291), .B(N239), .Z(n1397) );
  OR2 U2921 ( .A(n1396), .B(n1333), .Z(N833) );
  OR2 U2922 ( .A(n1394), .B(n1395), .Z(n1396) );
  OR2 U2923 ( .A(n1392), .B(n1393), .Z(n1395) );
  OR2 U2924 ( .A(n1390), .B(n1391), .Z(n1394) );
  OR2 U2925 ( .A(n1388), .B(n1389), .Z(n1393) );
  OR2 U2926 ( .A(n1386), .B(n1387), .Z(n1392) );
  OR2 U2927 ( .A(n1384), .B(n1385), .Z(n1391) );
  OR2 U2928 ( .A(n1382), .B(n1383), .Z(n1390) );
  OR2 U2929 ( .A(n1380), .B(n1381), .Z(n1389) );
  OR2 U2930 ( .A(n1378), .B(n1379), .Z(n1388) );
  OR2 U2931 ( .A(n1376), .B(n1377), .Z(n1387) );
  OR2 U2932 ( .A(n1374), .B(n1375), .Z(n1386) );
  OR2 U2933 ( .A(n1372), .B(n1373), .Z(n1385) );
  OR2 U2934 ( .A(n1370), .B(n1371), .Z(n1384) );
  OR2 U2935 ( .A(n1368), .B(n1369), .Z(n1383) );
  OR2 U2936 ( .A(n1366), .B(n1367), .Z(n1382) );
  OR2 U2937 ( .A(n1364), .B(n1365), .Z(n1381) );
  OR2 U2938 ( .A(n1362), .B(n1363), .Z(n1380) );
  OR2 U2939 ( .A(n1360), .B(n1361), .Z(n1379) );
  OR2 U2940 ( .A(n1358), .B(n1359), .Z(n1378) );
  OR2 U2941 ( .A(n1356), .B(n1357), .Z(n1377) );
  OR2 U2942 ( .A(n1354), .B(n1355), .Z(n1376) );
  OR2 U2943 ( .A(n1352), .B(n1353), .Z(n1375) );
  OR2 U2944 ( .A(n1350), .B(n1351), .Z(n1374) );
  OR2 U2945 ( .A(n1348), .B(n1349), .Z(n1373) );
  OR2 U2946 ( .A(n1346), .B(n1347), .Z(n1372) );
  OR2 U2947 ( .A(n1344), .B(n1345), .Z(n1371) );
  OR2 U2948 ( .A(n1342), .B(n1343), .Z(n1370) );
  OR2 U2949 ( .A(n1340), .B(n1341), .Z(n1369) );
  OR2 U2950 ( .A(n1338), .B(n1339), .Z(n1368) );
  OR2 U2951 ( .A(n1336), .B(n1337), .Z(n1367) );
  OR2 U2952 ( .A(n1334), .B(n1335), .Z(n1366) );
  OR2 U2953 ( .A(n1331), .B(n1332), .Z(n1365) );
  OR2 U2954 ( .A(n1329), .B(n1330), .Z(n1364) );
  OR2 U2955 ( .A(n1327), .B(n1328), .Z(n1363) );
  OR2 U2956 ( .A(n1325), .B(n1326), .Z(n1362) );
  OR2 U2957 ( .A(n1323), .B(n1324), .Z(n1361) );
  OR2 U2958 ( .A(n1321), .B(n1322), .Z(n1360) );
  OR2 U2959 ( .A(n1319), .B(n1320), .Z(n1359) );
  OR2 U2960 ( .A(n1317), .B(n1318), .Z(n1358) );
  OR2 U2961 ( .A(n1315), .B(n1316), .Z(n1357) );
  OR2 U2962 ( .A(n1313), .B(n1314), .Z(n1356) );
  OR2 U2963 ( .A(n1311), .B(n1312), .Z(n1355) );
  OR2 U2964 ( .A(n1309), .B(n1310), .Z(n1354) );
  OR2 U2965 ( .A(n1307), .B(n1308), .Z(n1353) );
  OR2 U2966 ( .A(n1305), .B(n1306), .Z(n1352) );
  OR2 U2967 ( .A(n1303), .B(n1304), .Z(n1351) );
  OR2 U2968 ( .A(n1301), .B(n1302), .Z(n1350) );
  OR2 U2969 ( .A(n1299), .B(n1300), .Z(n1349) );
  OR2 U2970 ( .A(n1297), .B(n1298), .Z(n1348) );
  OR2 U2971 ( .A(n1295), .B(n1296), .Z(n1347) );
  OR2 U2972 ( .A(n1293), .B(n1294), .Z(n1346) );
  OR2 U2973 ( .A(n1291), .B(n1292), .Z(n1345) );
  OR2 U2974 ( .A(n1289), .B(n1290), .Z(n1344) );
  OR2 U2975 ( .A(n1287), .B(n1288), .Z(n1343) );
  OR2 U2976 ( .A(n1174), .B(n1286), .Z(n1342) );
  OR2 U2977 ( .A(n1284), .B(n1285), .Z(n1341) );
  OR2 U2978 ( .A(n1282), .B(n1283), .Z(n1340) );
  OR2 U2979 ( .A(n1280), .B(n1281), .Z(n1339) );
  OR2 U2980 ( .A(n1278), .B(n1279), .Z(n1338) );
  OR2 U2981 ( .A(n1276), .B(n1277), .Z(n1337) );
  OR2 U2982 ( .A(n1274), .B(n1275), .Z(n1336) );
  OR2 U2983 ( .A(n1272), .B(n1273), .Z(n1335) );
  OR2 U2984 ( .A(n1270), .B(n1271), .Z(n1334) );
  OR2 U2985 ( .A(n1268), .B(n1269), .Z(n1333) );
  OR2 U2986 ( .A(n1266), .B(n1267), .Z(n1332) );
  OR2 U2987 ( .A(n1264), .B(n1265), .Z(n1331) );
  OR2 U2988 ( .A(n1262), .B(n1263), .Z(n1330) );
  OR2 U2989 ( .A(n1260), .B(n1261), .Z(n1329) );
  OR2 U2990 ( .A(n1258), .B(n1259), .Z(n1328) );
  OR2 U2991 ( .A(n1256), .B(n1257), .Z(n1327) );
  OR2 U2992 ( .A(n1254), .B(n1255), .Z(n1326) );
  OR2 U2993 ( .A(n1252), .B(n1253), .Z(n1325) );
  OR2 U2994 ( .A(n1250), .B(n1251), .Z(n1324) );
  OR2 U2995 ( .A(n1248), .B(n1249), .Z(n1323) );
  OR2 U2996 ( .A(n1246), .B(n1247), .Z(n1322) );
  OR2 U2997 ( .A(n1244), .B(n1245), .Z(n1321) );
  OR2 U2998 ( .A(n1242), .B(n1243), .Z(n1320) );
  OR2 U2999 ( .A(n1240), .B(n1241), .Z(n1319) );
  OR2 U3000 ( .A(n1238), .B(n1239), .Z(n1318) );
  OR2 U3001 ( .A(n1237), .B(N932), .Z(n1317) );
  OR2 U3002 ( .A(n1235), .B(n1236), .Z(n1316) );
  OR2 U3003 ( .A(n1233), .B(n1234), .Z(n1315) );
  OR2 U3004 ( .A(n1231), .B(n1232), .Z(n1314) );
  OR2 U3005 ( .A(n1229), .B(n1230), .Z(n1313) );
  OR2 U3006 ( .A(n1227), .B(n1228), .Z(n1312) );
  OR2 U3007 ( .A(n1225), .B(n1226), .Z(n1311) );
  OR2 U3008 ( .A(n1223), .B(n1224), .Z(n1310) );
  OR2 U3009 ( .A(n1221), .B(n1222), .Z(n1309) );
  OR2 U3010 ( .A(n1219), .B(n1220), .Z(n1308) );
  OR2 U3011 ( .A(n1217), .B(n1218), .Z(n1307) );
  OR2 U3012 ( .A(n1215), .B(n1216), .Z(n1306) );
  OR2 U3013 ( .A(n1213), .B(n1214), .Z(n1305) );
  OR2 U3014 ( .A(n1211), .B(n1212), .Z(n1304) );
  OR2 U3015 ( .A(n1209), .B(n1210), .Z(n1303) );
  OR2 U3016 ( .A(n1207), .B(n1208), .Z(n1302) );
  OR2 U3017 ( .A(n1205), .B(n1206), .Z(n1301) );
  OR2 U3018 ( .A(n1203), .B(n1204), .Z(n1300) );
  OR2 U3019 ( .A(n1201), .B(n1202), .Z(n1299) );
  OR2 U3020 ( .A(n1199), .B(n1200), .Z(n1298) );
  OR2 U3021 ( .A(n1197), .B(n1198), .Z(n1297) );
  OR2 U3022 ( .A(n1195), .B(n1196), .Z(n1296) );
  OR2 U3023 ( .A(n1193), .B(n1194), .Z(n1295) );
  OR2 U3024 ( .A(n1191), .B(n1192), .Z(n1294) );
  OR2 U3025 ( .A(n1189), .B(n1190), .Z(n1293) );
  OR2 U3026 ( .A(n1187), .B(n1188), .Z(n1292) );
  OR2 U3027 ( .A(n1185), .B(n1186), .Z(n1291) );
  OR2 U3028 ( .A(n1183), .B(n1184), .Z(n1290) );
  OR2 U3029 ( .A(n1181), .B(n1182), .Z(n1289) );
  OR2 U3030 ( .A(n1179), .B(n1180), .Z(n1288) );
  OR2 U3031 ( .A(n1177), .B(n1178), .Z(n1287) );
  OR2 U3032 ( .A(n1175), .B(n1176), .Z(n1286) );
  OR2 U3033 ( .A(n1172), .B(n1173), .Z(n1285) );
  OR2 U3034 ( .A(n1170), .B(n1171), .Z(n1284) );
  OR2 U3035 ( .A(n1168), .B(n1169), .Z(n1283) );
  OR2 U3036 ( .A(n1166), .B(n1167), .Z(n1282) );
  OR2 U3037 ( .A(n1164), .B(n1165), .Z(n1281) );
  OR2 U3038 ( .A(n1162), .B(n1163), .Z(n1280) );
  OR2 U3039 ( .A(n1160), .B(n1161), .Z(n1279) );
  OR2 U3040 ( .A(n1158), .B(n1159), .Z(n1278) );
  OR2 U3041 ( .A(n1156), .B(n1157), .Z(n1277) );
  OR2 U3042 ( .A(n1154), .B(n1155), .Z(n1276) );
  OR2 U3043 ( .A(n1152), .B(n1153), .Z(n1275) );
  OR2 U3044 ( .A(n1150), .B(n1151), .Z(n1274) );
  OR2 U3045 ( .A(n1148), .B(n1149), .Z(n1273) );
  OR2 U3046 ( .A(n1146), .B(n1147), .Z(n1272) );
  OR2 U3047 ( .A(n1144), .B(n1145), .Z(n1271) );
  OR2 U3048 ( .A(n1142), .B(n1143), .Z(n1270) );
  AN2 U3049 ( .A(pos_disp_tx), .B(N8311), .Z(n1269) );
  AN2 U3050 ( .A(pos_disp_tx), .B(n153), .Z(n1268) );
  AN2 U3051 ( .A(pos_disp_tx), .B(n33), .Z(n1267) );
  AN2 U3052 ( .A(n291), .B(n168), .Z(n1266) );
  AN2 U3053 ( .A(pos_disp_tx), .B(n19), .Z(n1265) );
  AN2 U3054 ( .A(n291), .B(n157), .Z(n1264) );
  AN2 U3055 ( .A(n291), .B(n37), .Z(n1263) );
  AN2 U3056 ( .A(pos_disp_tx), .B(n172), .Z(n1262) );
  AN2 U3057 ( .A(pos_disp_tx), .B(n26), .Z(n1261) );
  AN2 U3058 ( .A(n291), .B(n161), .Z(n1260) );
  AN2 U3059 ( .A(n291), .B(n40), .Z(n1259) );
  AN2 U3060 ( .A(n291), .B(n175), .Z(n1258) );
  AN2 U3061 ( .A(n291), .B(n30), .Z(n1257) );
  AN2 U3062 ( .A(n291), .B(n165), .Z(n1256) );
  AN2 U3063 ( .A(n291), .B(n43), .Z(n1255) );
  AN2 U3064 ( .A(pos_disp_tx), .B(n178), .Z(n1254) );
  AN2 U3065 ( .A(pos_disp_tx), .B(n23), .Z(n1253) );
  AN2 U3066 ( .A(n291), .B(n154), .Z(n1252) );
  AN2 U3067 ( .A(n291), .B(n34), .Z(n1251) );
  AN2 U3068 ( .A(n291), .B(n169), .Z(n1250) );
  AN2 U3069 ( .A(n291), .B(n20), .Z(n1249) );
  AN2 U3070 ( .A(n291), .B(n158), .Z(n1248) );
  AN2 U3071 ( .A(n291), .B(n38), .Z(n1247) );
  AN2 U3072 ( .A(pos_disp_tx), .B(n173), .Z(n1246) );
  AN2 U3073 ( .A(n291), .B(n27), .Z(n1245) );
  AN2 U3074 ( .A(n291), .B(n162), .Z(n1244) );
  AN2 U3075 ( .A(n291), .B(n41), .Z(n1243) );
  AN2 U3076 ( .A(pos_disp_tx), .B(n176), .Z(n1242) );
  AN2 U3077 ( .A(n291), .B(n31), .Z(n1241) );
  AN2 U3078 ( .A(pos_disp_tx), .B(n166), .Z(n1240) );
  AN2 U3079 ( .A(pos_disp_tx), .B(n44), .Z(n1239) );
  AN2 U3080 ( .A(pos_disp_tx), .B(n179), .Z(n1238) );
  AN2 U3081 ( .A(n291), .B(n62), .Z(n1237) );
  AN2 U3082 ( .A(n291), .B(n233), .Z(n1236) );
  AN2 U3083 ( .A(n291), .B(n99), .Z(n1235) );
  AN2 U3084 ( .A(pos_disp_tx), .B(n195), .Z(n1234) );
  AN2 U3085 ( .A(n291), .B(n50), .Z(n1233) );
  AN2 U3086 ( .A(pos_disp_tx), .B(n245), .Z(n1232) );
  AN2 U3087 ( .A(pos_disp_tx), .B(n111), .Z(n1231) );
  AN2 U3088 ( .A(n291), .B(n208), .Z(n1230) );
  AN2 U3089 ( .A(n291), .B(n74), .Z(n1229) );
  AN2 U3090 ( .A(pos_disp_tx), .B(n257), .Z(n1228) );
  AN2 U3091 ( .A(pos_disp_tx), .B(n123), .Z(n1227) );
  AN2 U3092 ( .A(pos_disp_tx), .B(n221), .Z(n1226) );
  AN2 U3093 ( .A(pos_disp_tx), .B(n87), .Z(n1225) );
  AN2 U3094 ( .A(pos_disp_tx), .B(n270), .Z(n1224) );
  AN2 U3095 ( .A(pos_disp_tx), .B(n136), .Z(n1223) );
  AN2 U3096 ( .A(n291), .B(n184), .Z(n1222) );
  AN2 U3097 ( .A(n291), .B(n63), .Z(n1221) );
  AN2 U3098 ( .A(pos_disp_tx), .B(n234), .Z(n1220) );
  AN2 U3099 ( .A(pos_disp_tx), .B(n100), .Z(n1219) );
  AN2 U3100 ( .A(pos_disp_tx), .B(n196), .Z(n1218) );
  AN2 U3101 ( .A(pos_disp_tx), .B(n51), .Z(n1217) );
  AN2 U3102 ( .A(pos_disp_tx), .B(n246), .Z(n1216) );
  AN2 U3103 ( .A(pos_disp_tx), .B(n112), .Z(n1215) );
  AN2 U3104 ( .A(n291), .B(n209), .Z(n1214) );
  AN2 U3105 ( .A(pos_disp_tx), .B(n75), .Z(n1213) );
  AN2 U3106 ( .A(pos_disp_tx), .B(n258), .Z(n1212) );
  AN2 U3107 ( .A(pos_disp_tx), .B(n124), .Z(n1211) );
  AN2 U3108 ( .A(n291), .B(n222), .Z(n1210) );
  AN2 U3109 ( .A(pos_disp_tx), .B(n88), .Z(n1209) );
  AN2 U3110 ( .A(n291), .B(n271), .Z(n1208) );
  AN2 U3111 ( .A(n291), .B(n137), .Z(n1207) );
  AN2 U3112 ( .A(n291), .B(n185), .Z(n1206) );
  AN2 U3113 ( .A(n291), .B(n64), .Z(n1205) );
  AN2 U3114 ( .A(n291), .B(n235), .Z(n1204) );
  AN2 U3115 ( .A(n291), .B(n101), .Z(n1203) );
  AN2 U3116 ( .A(pos_disp_tx), .B(n197), .Z(n1202) );
  AN2 U3117 ( .A(n291), .B(n52), .Z(n1201) );
  AN2 U3118 ( .A(pos_disp_tx), .B(n247), .Z(n1200) );
  AN2 U3119 ( .A(pos_disp_tx), .B(n113), .Z(n1199) );
  AN2 U3120 ( .A(n291), .B(n210), .Z(n1198) );
  AN2 U3121 ( .A(n291), .B(n76), .Z(n1197) );
  AN2 U3122 ( .A(pos_disp_tx), .B(n259), .Z(n1196) );
  AN2 U3123 ( .A(pos_disp_tx), .B(n125), .Z(n1195) );
  AN2 U3124 ( .A(pos_disp_tx), .B(n223), .Z(n1194) );
  AN2 U3125 ( .A(pos_disp_tx), .B(n89), .Z(n1193) );
  AN2 U3126 ( .A(pos_disp_tx), .B(n272), .Z(n1192) );
  AN2 U3127 ( .A(pos_disp_tx), .B(n138), .Z(n1191) );
  AN2 U3128 ( .A(n291), .B(n186), .Z(n1190) );
  AN2 U3129 ( .A(n291), .B(n65), .Z(n1189) );
  AN2 U3130 ( .A(pos_disp_tx), .B(n236), .Z(n1188) );
  AN2 U3131 ( .A(pos_disp_tx), .B(n102), .Z(n1187) );
  AN2 U3132 ( .A(pos_disp_tx), .B(n198), .Z(n1186) );
  AN2 U3133 ( .A(pos_disp_tx), .B(n53), .Z(n1185) );
  AN2 U3134 ( .A(pos_disp_tx), .B(n248), .Z(n1184) );
  AN2 U3135 ( .A(pos_disp_tx), .B(n114), .Z(n1183) );
  AN2 U3136 ( .A(n291), .B(n211), .Z(n1182) );
  AN2 U3137 ( .A(pos_disp_tx), .B(n77), .Z(n1181) );
  AN2 U3138 ( .A(pos_disp_tx), .B(n260), .Z(n1180) );
  AN2 U3139 ( .A(pos_disp_tx), .B(n126), .Z(n1179) );
  AN2 U3140 ( .A(n291), .B(n224), .Z(n1178) );
  AN2 U3141 ( .A(pos_disp_tx), .B(n90), .Z(n1177) );
  AN2 U3142 ( .A(n291), .B(n273), .Z(n1176) );
  AN2 U3143 ( .A(n291), .B(n139), .Z(n1175) );
  AN2 U3144 ( .A(n291), .B(n187), .Z(n1174) );
  AN2 U3145 ( .A(pos_disp_tx), .B(n70), .Z(n1173) );
  AN2 U3146 ( .A(pos_disp_tx), .B(n241), .Z(n1172) );
  AN2 U3147 ( .A(pos_disp_tx), .B(n107), .Z(n1171) );
  AN2 U3148 ( .A(n291), .B(n203), .Z(n1170) );
  AN2 U3149 ( .A(pos_disp_tx), .B(n58), .Z(n1169) );
  AN2 U3150 ( .A(n291), .B(n253), .Z(n1168) );
  AN2 U3151 ( .A(n291), .B(n119), .Z(n1167) );
  AN2 U3152 ( .A(pos_disp_tx), .B(n216), .Z(n1166) );
  AN2 U3153 ( .A(pos_disp_tx), .B(n82), .Z(n1165) );
  AN2 U3154 ( .A(n291), .B(n265), .Z(n1164) );
  AN2 U3155 ( .A(n291), .B(n131), .Z(n1163) );
  AN2 U3156 ( .A(n291), .B(n229), .Z(n1162) );
  AN2 U3157 ( .A(n291), .B(n95), .Z(n1161) );
  AN2 U3158 ( .A(n291), .B(n278), .Z(n1160) );
  AN2 U3159 ( .A(n291), .B(n144), .Z(n1159) );
  AN2 U3160 ( .A(pos_disp_tx), .B(n192), .Z(n1158) );
  AN2 U3161 ( .A(pos_disp_tx), .B(n71), .Z(n1157) );
  AN2 U3162 ( .A(n291), .B(n242), .Z(n1156) );
  AN2 U3163 ( .A(n291), .B(n108), .Z(n1155) );
  AN2 U3164 ( .A(n291), .B(n204), .Z(n1154) );
  AN2 U3165 ( .A(n291), .B(n59), .Z(n1153) );
  AN2 U3166 ( .A(n291), .B(n254), .Z(n1152) );
  AN2 U3167 ( .A(n291), .B(n120), .Z(n1151) );
  AN2 U3168 ( .A(pos_disp_tx), .B(n217), .Z(n1150) );
  AN2 U3169 ( .A(n291), .B(n83), .Z(n1149) );
  AN2 U3170 ( .A(n291), .B(n266), .Z(n1148) );
  AN2 U3171 ( .A(n291), .B(n132), .Z(n1147) );
  AN2 U3172 ( .A(pos_disp_tx), .B(n230), .Z(n1146) );
  AN2 U3173 ( .A(n291), .B(n96), .Z(n1145) );
  AN2 U3174 ( .A(pos_disp_tx), .B(n279), .Z(n1144) );
  AN2 U3175 ( .A(pos_disp_tx), .B(n145), .Z(n1143) );
  AN2 U3176 ( .A(pos_disp_tx), .B(N239), .Z(n1142) );
  OR2 U3177 ( .A(n1140), .B(n1141), .Z(N832) );
  OR2 U3178 ( .A(n1138), .B(n1139), .Z(n1141) );
  OR2 U3179 ( .A(n1136), .B(n1137), .Z(n1140) );
  OR2 U3180 ( .A(n1134), .B(n1135), .Z(n1139) );
  OR2 U3181 ( .A(n1132), .B(n1133), .Z(n1138) );
  OR2 U3182 ( .A(n1130), .B(n1131), .Z(n1137) );
  OR2 U3183 ( .A(n1128), .B(n1129), .Z(n1136) );
  OR2 U3184 ( .A(n1127), .B(n1112), .Z(n1135) );
  OR2 U3185 ( .A(n1125), .B(n1126), .Z(n1134) );
  OR2 U3186 ( .A(n1123), .B(n1124), .Z(n1133) );
  OR2 U3187 ( .A(n1121), .B(n1122), .Z(n1132) );
  OR2 U3188 ( .A(n1119), .B(n1120), .Z(n1131) );
  OR2 U3189 ( .A(n1117), .B(n1118), .Z(n1130) );
  OR2 U3190 ( .A(n1115), .B(n1116), .Z(n1129) );
  OR2 U3191 ( .A(n1113), .B(n1114), .Z(n1128) );
  OR2 U3192 ( .A(n1110), .B(n1111), .Z(n1127) );
  OR2 U3193 ( .A(n1108), .B(n1109), .Z(n1126) );
  OR2 U3194 ( .A(n1106), .B(n1107), .Z(n1125) );
  OR2 U3195 ( .A(n1104), .B(n1105), .Z(n1124) );
  OR2 U3196 ( .A(n1102), .B(n1103), .Z(n1123) );
  OR2 U3197 ( .A(n1100), .B(n1101), .Z(n1122) );
  OR2 U3198 ( .A(n1098), .B(n1099), .Z(n1121) );
  OR2 U3199 ( .A(n1096), .B(n1097), .Z(n1120) );
  OR2 U3200 ( .A(n1094), .B(n1095), .Z(n1119) );
  OR2 U3201 ( .A(n1092), .B(n1093), .Z(n1118) );
  OR2 U3202 ( .A(n1090), .B(n1091), .Z(n1117) );
  OR2 U3203 ( .A(n1088), .B(n1089), .Z(n1116) );
  OR2 U3204 ( .A(n1086), .B(n1087), .Z(n1115) );
  OR2 U3205 ( .A(n1084), .B(n1085), .Z(n1114) );
  OR2 U3206 ( .A(n1082), .B(n1083), .Z(n1113) );
  OR2 U3207 ( .A(n1080), .B(n1081), .Z(n1112) );
  OR2 U3208 ( .A(n1078), .B(n1079), .Z(n1111) );
  OR2 U3209 ( .A(n1076), .B(n1077), .Z(n1110) );
  OR2 U3210 ( .A(n1074), .B(n1075), .Z(n1109) );
  OR2 U3211 ( .A(n1072), .B(n1073), .Z(n1108) );
  OR2 U3212 ( .A(n1070), .B(n1071), .Z(n1107) );
  OR2 U3213 ( .A(n994), .B(n1069), .Z(n1106) );
  OR2 U3214 ( .A(n1067), .B(n1068), .Z(n1105) );
  OR2 U3215 ( .A(n1065), .B(n1066), .Z(n1104) );
  OR2 U3216 ( .A(n1063), .B(n1064), .Z(n1103) );
  OR2 U3217 ( .A(n1061), .B(n1062), .Z(n1102) );
  OR2 U3218 ( .A(n1059), .B(n1060), .Z(n1101) );
  OR2 U3219 ( .A(n1057), .B(n1058), .Z(n1100) );
  OR2 U3220 ( .A(n1055), .B(n1056), .Z(n1099) );
  OR2 U3221 ( .A(n1053), .B(n1054), .Z(n1098) );
  OR2 U3222 ( .A(n1051), .B(n1052), .Z(n1097) );
  OR2 U3223 ( .A(n1049), .B(n1050), .Z(n1096) );
  OR2 U3224 ( .A(n1047), .B(n1048), .Z(n1095) );
  OR2 U3225 ( .A(n1045), .B(n1046), .Z(n1094) );
  OR2 U3226 ( .A(n1043), .B(n1044), .Z(n1093) );
  OR2 U3227 ( .A(n1041), .B(n1042), .Z(n1092) );
  OR2 U3228 ( .A(n1039), .B(n1040), .Z(n1091) );
  OR2 U3229 ( .A(n1037), .B(n1038), .Z(n1090) );
  OR2 U3230 ( .A(n1035), .B(n1036), .Z(n1089) );
  OR2 U3231 ( .A(n1033), .B(n1034), .Z(n1088) );
  OR2 U3232 ( .A(n1031), .B(n1032), .Z(n1087) );
  OR2 U3233 ( .A(n1029), .B(n1030), .Z(n1086) );
  OR2 U3234 ( .A(n1027), .B(n1028), .Z(n1085) );
  OR2 U3235 ( .A(n1025), .B(n1026), .Z(n1084) );
  OR2 U3236 ( .A(n1023), .B(n1024), .Z(n1083) );
  OR2 U3237 ( .A(n1021), .B(n1022), .Z(n1082) );
  OR2 U3238 ( .A(n1019), .B(n1020), .Z(n1081) );
  OR2 U3239 ( .A(n1017), .B(n1018), .Z(n1080) );
  OR2 U3240 ( .A(n1015), .B(n1016), .Z(n1079) );
  OR2 U3241 ( .A(n1013), .B(n1014), .Z(n1078) );
  OR2 U3242 ( .A(n1011), .B(n1012), .Z(n1077) );
  OR2 U3243 ( .A(n1009), .B(n1010), .Z(n1076) );
  OR2 U3244 ( .A(n1007), .B(n1008), .Z(n1075) );
  OR2 U3245 ( .A(n1005), .B(n1006), .Z(n1074) );
  OR2 U3246 ( .A(n1003), .B(n1004), .Z(n1073) );
  OR2 U3247 ( .A(n1001), .B(n1002), .Z(n1072) );
  OR2 U3248 ( .A(n999), .B(n1000), .Z(n1071) );
  OR2 U3249 ( .A(n997), .B(n998), .Z(n1070) );
  OR2 U3250 ( .A(n995), .B(n996), .Z(n1069) );
  OR2 U3251 ( .A(n992), .B(n993), .Z(n1068) );
  OR2 U3252 ( .A(n990), .B(n991), .Z(n1067) );
  OR2 U3253 ( .A(n988), .B(n989), .Z(n1066) );
  OR2 U3254 ( .A(n986), .B(n987), .Z(n1065) );
  OR2 U3255 ( .A(n984), .B(n985), .Z(n1064) );
  OR2 U3256 ( .A(n982), .B(n983), .Z(n1063) );
  OR2 U3257 ( .A(n980), .B(n981), .Z(n1062) );
  OR2 U3258 ( .A(n978), .B(n979), .Z(n1061) );
  OR2 U3259 ( .A(n976), .B(n977), .Z(n1060) );
  OR2 U3260 ( .A(n974), .B(n975), .Z(n1059) );
  OR2 U3261 ( .A(n972), .B(n973), .Z(n1058) );
  OR2 U3262 ( .A(n970), .B(n971), .Z(n1057) );
  OR2 U3263 ( .A(n968), .B(n969), .Z(n1056) );
  OR2 U3264 ( .A(n966), .B(n967), .Z(n1055) );
  OR2 U3265 ( .A(n964), .B(n965), .Z(n1054) );
  OR2 U3266 ( .A(n962), .B(n963), .Z(n1053) );
  OR2 U3267 ( .A(n960), .B(n961), .Z(n1052) );
  OR2 U3268 ( .A(n958), .B(n959), .Z(n1051) );
  OR2 U3269 ( .A(n956), .B(n957), .Z(n1050) );
  OR2 U3270 ( .A(n954), .B(n955), .Z(n1049) );
  OR2 U3271 ( .A(n952), .B(n953), .Z(n1048) );
  OR2 U3272 ( .A(n950), .B(n951), .Z(n1047) );
  OR2 U3273 ( .A(n948), .B(n949), .Z(n1046) );
  OR2 U3274 ( .A(n946), .B(n947), .Z(n1045) );
  OR2 U3275 ( .A(n944), .B(n945), .Z(n1044) );
  OR2 U3276 ( .A(n942), .B(n943), .Z(n1043) );
  OR2 U3277 ( .A(n940), .B(n941), .Z(n1042) );
  OR2 U3278 ( .A(n938), .B(n939), .Z(n1041) );
  OR2 U3279 ( .A(n936), .B(n937), .Z(n1040) );
  OR2 U3280 ( .A(n934), .B(n935), .Z(n1039) );
  OR2 U3281 ( .A(n932), .B(n933), .Z(n1038) );
  OR2 U3282 ( .A(N908), .B(n931), .Z(n1037) );
  OR2 U3283 ( .A(n929), .B(n930), .Z(n1036) );
  OR2 U3284 ( .A(n927), .B(n928), .Z(n1035) );
  OR2 U3285 ( .A(n925), .B(n926), .Z(n1034) );
  OR2 U3286 ( .A(n923), .B(n924), .Z(n1033) );
  OR2 U3287 ( .A(n921), .B(n922), .Z(n1032) );
  OR2 U3288 ( .A(n919), .B(n920), .Z(n1031) );
  OR2 U3289 ( .A(n917), .B(n918), .Z(n1030) );
  OR2 U3290 ( .A(n915), .B(n916), .Z(n1029) );
  OR2 U3291 ( .A(n913), .B(n914), .Z(n1028) );
  OR2 U3292 ( .A(n911), .B(n912), .Z(n1027) );
  OR2 U3293 ( .A(n909), .B(n910), .Z(n1026) );
  OR2 U3294 ( .A(n907), .B(n908), .Z(n1025) );
  OR2 U3295 ( .A(n905), .B(n906), .Z(n1024) );
  OR2 U3296 ( .A(n903), .B(n904), .Z(n1023) );
  OR2 U3297 ( .A(n901), .B(n902), .Z(n1022) );
  OR2 U3298 ( .A(n899), .B(n900), .Z(n1021) );
  AN2 U3299 ( .A(n291), .B(N8311), .Z(n1020) );
  AN2 U3300 ( .A(n291), .B(n153), .Z(n1019) );
  AN2 U3301 ( .A(n291), .B(n33), .Z(n1018) );
  AN2 U3302 ( .A(pos_disp_tx), .B(n168), .Z(n1017) );
  AN2 U3303 ( .A(n291), .B(n19), .Z(n1016) );
  AN2 U3304 ( .A(pos_disp_tx), .B(n157), .Z(n1015) );
  AN2 U3305 ( .A(pos_disp_tx), .B(n37), .Z(n1014) );
  AN2 U3306 ( .A(n291), .B(n172), .Z(n1013) );
  AN2 U3307 ( .A(n291), .B(n26), .Z(n1012) );
  AN2 U3308 ( .A(pos_disp_tx), .B(n161), .Z(n1011) );
  AN2 U3309 ( .A(pos_disp_tx), .B(n40), .Z(n1010) );
  AN2 U3310 ( .A(pos_disp_tx), .B(n30), .Z(n1009) );
  AN2 U3311 ( .A(n291), .B(n178), .Z(n1008) );
  AN2 U3312 ( .A(n291), .B(n23), .Z(n1007) );
  AN2 U3313 ( .A(pos_disp_tx), .B(n169), .Z(n1006) );
  AN2 U3314 ( .A(pos_disp_tx), .B(n158), .Z(n1005) );
  AN2 U3315 ( .A(pos_disp_tx), .B(n38), .Z(n1004) );
  AN2 U3316 ( .A(n291), .B(n173), .Z(n1003) );
  AN2 U3317 ( .A(pos_disp_tx), .B(n27), .Z(n1002) );
  AN2 U3318 ( .A(pos_disp_tx), .B(n162), .Z(n1001) );
  AN2 U3319 ( .A(pos_disp_tx), .B(n41), .Z(n1000) );
  AN2 U3320 ( .A(n291), .B(n176), .Z(n999) );
  AN2 U3321 ( .A(pos_disp_tx), .B(n31), .Z(n998) );
  AN2 U3322 ( .A(n291), .B(n166), .Z(n997) );
  AN2 U3323 ( .A(n291), .B(n44), .Z(n996) );
  AN2 U3324 ( .A(n291), .B(n179), .Z(n995) );
  AN2 U3325 ( .A(pos_disp_tx), .B(n62), .Z(n994) );
  AN2 U3326 ( .A(pos_disp_tx), .B(n233), .Z(n993) );
  AN2 U3327 ( .A(pos_disp_tx), .B(n99), .Z(n992) );
  AN2 U3328 ( .A(n291), .B(n195), .Z(n991) );
  AN2 U3329 ( .A(pos_disp_tx), .B(n50), .Z(n990) );
  AN2 U3330 ( .A(n291), .B(n245), .Z(n989) );
  AN2 U3331 ( .A(n291), .B(n111), .Z(n988) );
  AN2 U3332 ( .A(pos_disp_tx), .B(n208), .Z(n987) );
  AN2 U3333 ( .A(pos_disp_tx), .B(n74), .Z(n986) );
  AN2 U3334 ( .A(n291), .B(n257), .Z(n985) );
  AN2 U3335 ( .A(n291), .B(n123), .Z(n984) );
  AN2 U3336 ( .A(n291), .B(n221), .Z(n983) );
  AN2 U3337 ( .A(n291), .B(n87), .Z(n982) );
  AN2 U3338 ( .A(n291), .B(n270), .Z(n981) );
  AN2 U3339 ( .A(n291), .B(n136), .Z(n980) );
  AN2 U3340 ( .A(pos_disp_tx), .B(n184), .Z(n979) );
  AN2 U3341 ( .A(pos_disp_tx), .B(n63), .Z(n978) );
  AN2 U3342 ( .A(n291), .B(n234), .Z(n977) );
  AN2 U3343 ( .A(n291), .B(n100), .Z(n976) );
  AN2 U3344 ( .A(n291), .B(n196), .Z(n975) );
  AN2 U3345 ( .A(n291), .B(n51), .Z(n974) );
  AN2 U3346 ( .A(n291), .B(n246), .Z(n973) );
  AN2 U3347 ( .A(n291), .B(n112), .Z(n972) );
  AN2 U3348 ( .A(pos_disp_tx), .B(n209), .Z(n971) );
  AN2 U3349 ( .A(n291), .B(n75), .Z(n970) );
  AN2 U3350 ( .A(n291), .B(n258), .Z(n969) );
  AN2 U3351 ( .A(n291), .B(n124), .Z(n968) );
  AN2 U3352 ( .A(pos_disp_tx), .B(n222), .Z(n967) );
  AN2 U3353 ( .A(n291), .B(n88), .Z(n966) );
  AN2 U3354 ( .A(pos_disp_tx), .B(n271), .Z(n965) );
  AN2 U3355 ( .A(pos_disp_tx), .B(n137), .Z(n964) );
  AN2 U3356 ( .A(pos_disp_tx), .B(n185), .Z(n963) );
  AN2 U3357 ( .A(n291), .B(n64), .Z(n962) );
  AN2 U3358 ( .A(n291), .B(n235), .Z(n961) );
  AN2 U3359 ( .A(n291), .B(n101), .Z(n960) );
  AN2 U3360 ( .A(pos_disp_tx), .B(n197), .Z(n959) );
  AN2 U3361 ( .A(n291), .B(n52), .Z(n958) );
  AN2 U3362 ( .A(pos_disp_tx), .B(n247), .Z(n957) );
  AN2 U3363 ( .A(pos_disp_tx), .B(n113), .Z(n956) );
  AN2 U3364 ( .A(n291), .B(n210), .Z(n955) );
  AN2 U3365 ( .A(n291), .B(n76), .Z(n954) );
  AN2 U3366 ( .A(pos_disp_tx), .B(n259), .Z(n953) );
  AN2 U3367 ( .A(pos_disp_tx), .B(n125), .Z(n952) );
  AN2 U3368 ( .A(pos_disp_tx), .B(n223), .Z(n951) );
  AN2 U3369 ( .A(pos_disp_tx), .B(n89), .Z(n950) );
  AN2 U3370 ( .A(pos_disp_tx), .B(n272), .Z(n949) );
  AN2 U3371 ( .A(pos_disp_tx), .B(n138), .Z(n948) );
  AN2 U3372 ( .A(n291), .B(n186), .Z(n947) );
  AN2 U3373 ( .A(n291), .B(n65), .Z(n946) );
  AN2 U3374 ( .A(pos_disp_tx), .B(n236), .Z(n945) );
  AN2 U3375 ( .A(pos_disp_tx), .B(n102), .Z(n944) );
  AN2 U3376 ( .A(pos_disp_tx), .B(n198), .Z(n943) );
  AN2 U3377 ( .A(pos_disp_tx), .B(n53), .Z(n942) );
  AN2 U3378 ( .A(pos_disp_tx), .B(n248), .Z(n941) );
  AN2 U3379 ( .A(pos_disp_tx), .B(n114), .Z(n940) );
  AN2 U3380 ( .A(n291), .B(n211), .Z(n939) );
  AN2 U3381 ( .A(pos_disp_tx), .B(n77), .Z(n938) );
  AN2 U3382 ( .A(pos_disp_tx), .B(n260), .Z(n937) );
  AN2 U3383 ( .A(pos_disp_tx), .B(n126), .Z(n936) );
  AN2 U3384 ( .A(n291), .B(n224), .Z(n935) );
  AN2 U3385 ( .A(pos_disp_tx), .B(n90), .Z(n934) );
  AN2 U3386 ( .A(n291), .B(n273), .Z(n933) );
  AN2 U3387 ( .A(n291), .B(n139), .Z(n932) );
  AN2 U3388 ( .A(n291), .B(n187), .Z(n931) );
  AN2 U3389 ( .A(pos_disp_tx), .B(n70), .Z(n930) );
  AN2 U3390 ( .A(pos_disp_tx), .B(n241), .Z(n929) );
  AN2 U3391 ( .A(pos_disp_tx), .B(n107), .Z(n928) );
  AN2 U3392 ( .A(n291), .B(n203), .Z(n927) );
  AN2 U3393 ( .A(pos_disp_tx), .B(n58), .Z(n926) );
  AN2 U3394 ( .A(n291), .B(n253), .Z(n925) );
  AN2 U3395 ( .A(n291), .B(n119), .Z(n924) );
  AN2 U3396 ( .A(pos_disp_tx), .B(n216), .Z(n923) );
  AN2 U3397 ( .A(pos_disp_tx), .B(n82), .Z(n922) );
  AN2 U3398 ( .A(n291), .B(n265), .Z(n921) );
  AN2 U3399 ( .A(n291), .B(n131), .Z(n920) );
  AN2 U3400 ( .A(n291), .B(n229), .Z(n919) );
  AN2 U3401 ( .A(n291), .B(n95), .Z(n918) );
  AN2 U3402 ( .A(n291), .B(n278), .Z(n917) );
  AN2 U3403 ( .A(n291), .B(n144), .Z(n916) );
  AN2 U3404 ( .A(pos_disp_tx), .B(n192), .Z(n915) );
  AN2 U3405 ( .A(pos_disp_tx), .B(n71), .Z(n914) );
  AN2 U3406 ( .A(n291), .B(n242), .Z(n913) );
  AN2 U3407 ( .A(n291), .B(n108), .Z(n912) );
  AN2 U3408 ( .A(n291), .B(n204), .Z(n911) );
  AN2 U3409 ( .A(n291), .B(n59), .Z(n910) );
  AN2 U3410 ( .A(n291), .B(n254), .Z(n909) );
  AN2 U3411 ( .A(n291), .B(n120), .Z(n908) );
  AN2 U3412 ( .A(pos_disp_tx), .B(n217), .Z(n907) );
  AN2 U3413 ( .A(n291), .B(n83), .Z(n906) );
  AN2 U3414 ( .A(n291), .B(n266), .Z(n905) );
  AN2 U3415 ( .A(n291), .B(n132), .Z(n904) );
  AN2 U3416 ( .A(pos_disp_tx), .B(n230), .Z(n903) );
  AN2 U3417 ( .A(n291), .B(n96), .Z(n902) );
  AN2 U3418 ( .A(pos_disp_tx), .B(n279), .Z(n901) );
  AN2 U3419 ( .A(pos_disp_tx), .B(n145), .Z(n900) );
  AN2 U3420 ( .A(pos_disp_tx), .B(N239), .Z(n899) );
  AN2 U3421 ( .A(N6341), .B(n290), .Z(pos_disp_tx_p) );
  OR2 U3422 ( .A(n896), .B(n897), .Z(N6341) );
  AN2 U3423 ( .A(N6331), .B(special_enc_in), .Z(n897) );
  AN2 U3424 ( .A(N6231), .B(n304), .Z(n896) );
  OR2 U3425 ( .A(n894), .B(n895), .Z(N6331) );
  AN2 U3426 ( .A(pos_disp_tx), .B(N6371), .Z(n895) );
  AN2 U3427 ( .A(n291), .B(N6351), .Z(n894) );
  OR2 U3428 ( .A(n892), .B(n893), .Z(N6231) );
  AN2 U3429 ( .A(n291), .B(n147), .Z(n893) );
  AN2 U3430 ( .A(pos_disp_tx), .B(N6721), .Z(n892) );
  AN2 U3431 ( .A(pos_disp_tx_p), .B(N2103), .Z(n891) );
  OR2 U3432 ( .A(n889), .B(n307), .Z(n890) );
  AN2 U3433 ( .A(tx_10bdata_todiag[9]), .B(N5103), .Z(n889) );
  AN2 U3434 ( .A(tx_10bdata_todiag[8]), .B(N5103), .Z(n888) );
  OR2 U3435 ( .A(n887), .B(N1190), .Z(tx_10bdata_predel[7]) );
  OR2 U3436 ( .A(n886), .B(n307), .Z(n887) );
  AN2 U3437 ( .A(tx_10bdata_todiag[7]), .B(N5103), .Z(n886) );
  OR2 U3438 ( .A(n885), .B(N1190), .Z(tx_10bdata_predel[6]) );
  AN2 U3439 ( .A(tx_10bdata_todiag[6]), .B(N5103), .Z(n885) );
  OR2 U3440 ( .A(n884), .B(N1190), .Z(tx_10bdata_predel[5]) );
  OR2 U3441 ( .A(n883), .B(n307), .Z(n884) );
  AN2 U3442 ( .A(tx_10bdata_todiag[5]), .B(N5103), .Z(n883) );
  OR2 U3443 ( .A(n882), .B(N1190), .Z(tx_10bdata_predel[4]) );
  AN2 U3444 ( .A(tx_10bdata_todiag[4]), .B(N5103), .Z(n882) );
  OR2 U3445 ( .A(n881), .B(N1190), .Z(tx_10bdata_predel[3]) );
  OR2 U3446 ( .A(n880), .B(n307), .Z(n881) );
  AN2 U3447 ( .A(tx_10bdata_todiag[3]), .B(N5103), .Z(n880) );
  AN2 U3448 ( .A(tx_10bdata_todiag[2]), .B(N5103), .Z(n879) );
  OR2 U3449 ( .A(n877), .B(n307), .Z(n878) );
  AN2 U3450 ( .A(tx_10bdata_todiag[1]), .B(N5103), .Z(n877) );
  AN2 U3451 ( .A(tx_10bdata_todiag[0]), .B(N5103), .Z(n876) );
  OR2 U3452 ( .A(n874), .B(n875), .Z(tx_enc_sel[3]) );
  AN2 U3453 ( .A(tx_enc_ctrl_sel_reg[3]), .B(link_up_loc), .Z(n875) );
  AN2 U3454 ( .A(tx_enc_conf_sel[3]), .B(N2105), .Z(n874) );
  OR2 U3455 ( .A(n872), .B(n873), .Z(tx_enc_sel[2]) );
  AN2 U3456 ( .A(tx_enc_ctrl_sel_reg[2]), .B(link_up_loc), .Z(n873) );
  AN2 U3457 ( .A(tx_enc_conf_sel[2]), .B(N2105), .Z(n872) );
  OR2 U3458 ( .A(n870), .B(n871), .Z(tx_enc_sel[1]) );
  AN2 U3459 ( .A(tx_enc_ctrl_sel_reg[1]), .B(link_up_loc), .Z(n871) );
  AN2 U3460 ( .A(tx_enc_conf_sel[1]), .B(N2105), .Z(n870) );
  OR2 U3461 ( .A(n868), .B(n869), .Z(tx_enc_sel[0]) );
  AN2 U3462 ( .A(tx_enc_ctrl_sel_reg[0]), .B(link_up_loc), .Z(n869) );
  AN2 U3463 ( .A(tx_enc_conf_sel[0]), .B(N2105), .Z(n868) );
  IV U3465 ( .A(N593), .Z(n99) );
  IV U3466 ( .A(N80), .Z(n9) );
  IV U3467 ( .A(N268), .Z(n83) );
  IV U3468 ( .A(N3101), .Z(n82) );
  IV U3469 ( .A(N73), .Z(n8) );
  IV U3470 ( .A(N480), .Z(n77) );
  IV U3471 ( .A(N514), .Z(n76) );
  IV U3472 ( .A(N548), .Z(n75) );
  IV U3473 ( .A(N5811), .Z(n74) );
  IV U3474 ( .A(N2911), .Z(n71) );
  IV U3475 ( .A(N329), .Z(n70) );
  IV U3476 ( .A(N67), .Z(n7) );
  IV U3477 ( .A(N496), .Z(n65) );
  IV U3478 ( .A(N530), .Z(n64) );
  IV U3479 ( .A(N564), .Z(n63) );
  IV U3480 ( .A(N597), .Z(n62) );
  IV U3481 ( .A(N62), .Z(n6) );
  IV U3482 ( .A(N319), .Z(n58) );
  IV U3483 ( .A(N522), .Z(n52) );
  IV U3484 ( .A(N589), .Z(n50) );
  IV U3485 ( .A(N57), .Z(n5) );
  IV U3486 ( .A(N7411), .Z(n44) );
  IV U3487 ( .A(N52), .Z(n4) );
  IV U3488 ( .A(N820), .Z(n33) );
  IV U3489 ( .A(jitter_study_tx[0]), .Z(n308) );
  IV U3490 ( .A(N6103), .Z(n307) );
  IV U3491 ( .A(jitter_study_tx[1]), .Z(n306) );
  IV U3492 ( .A(N8102), .Z(n305) );
  IV U3493 ( .A(special_enc_in), .Z(n304) );
  IV U3494 ( .A(encoder_sel[3]), .Z(n303) );
  IV U3495 ( .A(encoder_sel[2]), .Z(n302) );
  IV U3496 ( .A(encoder_sel[1]), .Z(n301) );
  IV U3497 ( .A(N848), .Z(n300) );
  IV U3498 ( .A(tx_enc_sel[3]), .Z(n3) );
  IV U3499 ( .A(N850), .Z(n298) );
  IV U3500 ( .A(N864), .Z(n297) );
  IV U3501 ( .A(encoder_sel[0]), .Z(n296) );
  IV U3502 ( .A(N8611), .Z(n295) );
  IV U3503 ( .A(N852), .Z(n293) );
  IV U3504 ( .A(pos_disp_tx), .Z(n291) );
  IV U3505 ( .A(rst_reg), .Z(n290) );
  IV U3506 ( .A(tx_8b_enc_in[7]), .Z(n289) );
  IV U3507 ( .A(tx_8b_enc_in[6]), .Z(n288) );
  IV U3508 ( .A(tx_8b_enc_in[5]), .Z(n287) );
  IV U3509 ( .A(tx_8b_enc_in[4]), .Z(n286) );
  IV U3510 ( .A(tx_8b_enc_in[3]), .Z(n285) );
  IV U3511 ( .A(tx_8b_enc_in[2]), .Z(n284) );
  IV U3512 ( .A(tx_8b_enc_in[1]), .Z(n283) );
  IV U3513 ( .A(N6061), .Z(n282) );
  IV U3514 ( .A(N6012), .Z(n281) );
  IV U3515 ( .A(N250), .Z(n279) );
  IV U3516 ( .A(N470), .Z(n273) );
  IV U3517 ( .A(N538), .Z(n271) );
  IV U3518 ( .A(N765), .Z(n27) );
  IV U3519 ( .A(N806), .Z(n26) );
  IV U3520 ( .A(N327), .Z(n241) );
  IV U3521 ( .A(N528), .Z(n235) );
  IV U3522 ( .A(N595), .Z(n233) );
  IV U3523 ( .A(N258), .Z(n230) );
  IV U3524 ( .A(N788), .Z(n23) );
  IV U3525 ( .A(N474), .Z(n224) );
  IV U3526 ( .A(N542), .Z(n222) );
  IV U3527 ( .A(N272), .Z(n217) );
  IV U3528 ( .A(N3121), .Z(n216) );
  IV U3529 ( .A(N482), .Z(n211) );
  IV U3530 ( .A(N516), .Z(n210) );
  IV U3531 ( .A(N550), .Z(n209) );
  IV U3532 ( .A(N583), .Z(n208) );
  IV U3533 ( .A(N97), .Z(n2) );
  IV U3534 ( .A(N296), .Z(n192) );
  IV U3535 ( .A(N815), .Z(n19) );
  IV U3536 ( .A(N466), .Z(n187) );
  IV U3537 ( .A(N500), .Z(n186) );
  IV U3538 ( .A(N534), .Z(n185) );
  IV U3539 ( .A(N567), .Z(n184) );
  IV U3540 ( .A(txd_d[3]), .Z(n18) );
  IV U3541 ( .A(N737), .Z(n179) );
  IV U3542 ( .A(N792), .Z(n178) );
  IV U3543 ( .A(N755), .Z(n176) );
  IV U3544 ( .A(N769), .Z(n173) );
  IV U3545 ( .A(N808), .Z(n172) );
  IV U3546 ( .A(txd_d[2]), .Z(n17) );
  IV U3547 ( .A(N817), .Z(n168) );
  IV U3548 ( .A(N748), .Z(n166) );
  IV U3549 ( .A(txd_d[1]), .Z(n16) );
  IV U3550 ( .A(N8121), .Z(n157) );
  IV U3551 ( .A(N823), .Z(n153) );
  IV U3552 ( .A(tx_8b_enc_in[0]), .Z(n152) );
  IV U3553 ( .A(n3407), .Z(n150) );
  AN2 U3554 ( .A(n3408), .B(n3409), .Z(n3407) );
  AN2 U3555 ( .A(n3410), .B(N5761), .Z(n3409) );
  AN2 U3556 ( .A(N5701), .B(N5501), .Z(n3410) );
  AN2 U3557 ( .A(N5971), .B(N5951), .Z(n3408) );
  IV U3558 ( .A(txd_d[0]), .Z(n15) );
  IV U3559 ( .A(n3411), .Z(n148) );
  AN2 U3560 ( .A(n3412), .B(n3413), .Z(n3411) );
  AN2 U3561 ( .A(n3414), .B(n3415), .Z(n3413) );
  AN2 U3562 ( .A(n3416), .B(n3417), .Z(n3415) );
  AN2 U3563 ( .A(n3418), .B(n3419), .Z(n3417) );
  AN2 U3564 ( .A(n3420), .B(n3421), .Z(n3419) );
  AN2 U3565 ( .A(n3422), .B(n3423), .Z(n3421) );
  AN2 U3566 ( .A(N10110), .B(n3424), .Z(n3423) );
  IV U3567 ( .A(N3010), .Z(n3424) );
  AN2 U3568 ( .A(N11110), .B(N10710), .Z(n3422) );
  AN2 U3569 ( .A(n3425), .B(n3426), .Z(n3420) );
  AN2 U3570 ( .A(N11510), .B(N11310), .Z(n3426) );
  AN2 U3571 ( .A(N1291), .B(N1251), .Z(n3425) );
  AN2 U3572 ( .A(n3427), .B(n3428), .Z(n3418) );
  AN2 U3573 ( .A(n3429), .B(n3430), .Z(n3428) );
  AN2 U3574 ( .A(N1331), .B(N1312), .Z(n3430) );
  AN2 U3575 ( .A(N1401), .B(N1381), .Z(n3429) );
  AN2 U3576 ( .A(n3431), .B(n3432), .Z(n3427) );
  AN2 U3577 ( .A(N1441), .B(N1421), .Z(n3432) );
  AN2 U3578 ( .A(N1481), .B(N1461), .Z(n3431) );
  AN2 U3579 ( .A(n3433), .B(n3434), .Z(n3416) );
  AN2 U3580 ( .A(n3435), .B(n3436), .Z(n3434) );
  AN2 U3581 ( .A(n3437), .B(n3438), .Z(n3436) );
  AN2 U3582 ( .A(N1591), .B(N1571), .Z(n3438) );
  AN2 U3583 ( .A(N1631), .B(N1612), .Z(n3437) );
  AN2 U3584 ( .A(n3439), .B(n3440), .Z(n3435) );
  AN2 U3585 ( .A(N1671), .B(N1651), .Z(n3440) );
  AN2 U3586 ( .A(N1751), .B(N1731), .Z(n3439) );
  AN2 U3587 ( .A(n3441), .B(n3442), .Z(n3433) );
  AN2 U3588 ( .A(n3443), .B(n3444), .Z(n3442) );
  AN2 U3589 ( .A(N1951), .B(N1791), .Z(n3444) );
  AN2 U3590 ( .A(N2012), .B(N1991), .Z(n3443) );
  AN2 U3591 ( .A(n3445), .B(n3446), .Z(n3441) );
  AN2 U3592 ( .A(N2071), .B(N2031), .Z(n3446) );
  AN2 U3593 ( .A(N2112), .B(N2091), .Z(n3445) );
  AN2 U3594 ( .A(n3447), .B(n3448), .Z(n3414) );
  AN2 U3595 ( .A(n3449), .B(n3450), .Z(n3448) );
  AN2 U3596 ( .A(n3451), .B(n3452), .Z(n3450) );
  AN2 U3597 ( .A(n3453), .B(n3454), .Z(n3452) );
  AN2 U3598 ( .A(N2152), .B(N2132), .Z(n3454) );
  AN2 U3599 ( .A(N2241), .B(N2171), .Z(n3453) );
  AN2 U3600 ( .A(n3455), .B(n3456), .Z(n3451) );
  AN2 U3601 ( .A(N2281), .B(N2261), .Z(n3456) );
  AN2 U3602 ( .A(N2321), .B(N2301), .Z(n3455) );
  AN2 U3603 ( .A(n3457), .B(n3458), .Z(n3449) );
  AN2 U3604 ( .A(n3459), .B(n3460), .Z(n3458) );
  AN2 U3605 ( .A(N2401), .B(N2341), .Z(n3460) );
  AN2 U3606 ( .A(N2461), .B(N2421), .Z(n3459) );
  AN2 U3607 ( .A(n3461), .B(n3462), .Z(n3457) );
  AN2 U3608 ( .A(N2651), .B(N2612), .Z(n3462) );
  AN2 U3609 ( .A(N2691), .B(N2671), .Z(n3461) );
  AN2 U3610 ( .A(n3463), .B(n3464), .Z(n3447) );
  AN2 U3611 ( .A(n3465), .B(n3466), .Z(n3464) );
  AN2 U3612 ( .A(n3467), .B(n3468), .Z(n3466) );
  AN2 U3613 ( .A(N2751), .B(N2731), .Z(n3468) );
  AN2 U3614 ( .A(N2791), .B(N2771), .Z(n3467) );
  AN2 U3615 ( .A(n3469), .B(n3470), .Z(n3465) );
  AN2 U3616 ( .A(N2831), .B(N2812), .Z(n3470) );
  AN2 U3617 ( .A(N2921), .B(N2901), .Z(n3469) );
  AN2 U3618 ( .A(n3471), .B(n3472), .Z(n3463) );
  AN2 U3619 ( .A(n3473), .B(n3474), .Z(n3472) );
  AN2 U3620 ( .A(N2961), .B(N2941), .Z(n3474) );
  AN2 U3621 ( .A(N3001), .B(N2981), .Z(n3473) );
  AN2 U3622 ( .A(n3475), .B(N3110), .Z(n3471) );
  AN2 U3623 ( .A(N3081), .B(N3061), .Z(n3475) );
  AN2 U3624 ( .A(n3476), .B(n3477), .Z(n3412) );
  AN2 U3625 ( .A(n3478), .B(n3479), .Z(n3477) );
  AN2 U3626 ( .A(n3480), .B(n3481), .Z(n3479) );
  AN2 U3627 ( .A(n3482), .B(n3483), .Z(n3481) );
  AN2 U3628 ( .A(n3484), .B(n3485), .Z(n3483) );
  AN2 U3629 ( .A(N3201), .B(N3122), .Z(n3485) );
  AN2 U3630 ( .A(N3241), .B(N3221), .Z(n3484) );
  AN2 U3631 ( .A(n3486), .B(n3487), .Z(n3482) );
  AN2 U3632 ( .A(N3310), .B(N3301), .Z(n3487) );
  AN2 U3633 ( .A(N3521), .B(N3381), .Z(n3486) );
  AN2 U3634 ( .A(n3488), .B(n3489), .Z(n3480) );
  AN2 U3635 ( .A(n3490), .B(n3491), .Z(n3489) );
  AN2 U3636 ( .A(N3691), .B(N3541), .Z(n3491) );
  AN2 U3637 ( .A(N3771), .B(N3712), .Z(n3490) );
  AN2 U3638 ( .A(n3492), .B(n3493), .Z(n3488) );
  AN2 U3639 ( .A(N3831), .B(N3812), .Z(n3493) );
  AN2 U3640 ( .A(N3941), .B(N3851), .Z(n3492) );
  AN2 U3641 ( .A(n3494), .B(n3495), .Z(n3478) );
  AN2 U3642 ( .A(n3496), .B(n3497), .Z(n3495) );
  AN2 U3643 ( .A(n3498), .B(n3499), .Z(n3497) );
  AN2 U3644 ( .A(N4001), .B(N3981), .Z(n3499) );
  AN2 U3645 ( .A(N4061), .B(N4021), .Z(n3498) );
  AN2 U3646 ( .A(n3500), .B(n3501), .Z(n3496) );
  AN2 U3647 ( .A(N4102), .B(N4081), .Z(n3501) );
  AN2 U3648 ( .A(N4141), .B(N4122), .Z(n3500) );
  AN2 U3649 ( .A(n3502), .B(n3503), .Z(n3494) );
  AN2 U3650 ( .A(n3504), .B(n3505), .Z(n3503) );
  AN2 U3651 ( .A(N4210), .B(N4161), .Z(n3505) );
  AN2 U3652 ( .A(N4251), .B(N4231), .Z(n3504) );
  AN2 U3653 ( .A(n3506), .B(N4312), .Z(n3502) );
  AN2 U3654 ( .A(N4291), .B(N4271), .Z(n3506) );
  AN2 U3655 ( .A(n3507), .B(n3508), .Z(n3476) );
  AN2 U3656 ( .A(n3509), .B(n3510), .Z(n3508) );
  AN2 U3657 ( .A(n3511), .B(n3512), .Z(n3510) );
  AN2 U3658 ( .A(n3513), .B(n3514), .Z(n3512) );
  AN2 U3659 ( .A(N4391), .B(N4331), .Z(n3514) );
  AN2 U3660 ( .A(N4451), .B(N4412), .Z(n3513) );
  AN2 U3661 ( .A(n3515), .B(n3516), .Z(n3511) );
  AN2 U3662 ( .A(N4661), .B(N4612), .Z(n3516) );
  AN2 U3663 ( .A(N4701), .B(N4681), .Z(n3515) );
  AN2 U3664 ( .A(n3517), .B(n3518), .Z(n3509) );
  AN2 U3665 ( .A(n3519), .B(n3520), .Z(n3518) );
  AN2 U3666 ( .A(N4771), .B(N4751), .Z(n3520) );
  AN2 U3667 ( .A(N4812), .B(N4791), .Z(n3519) );
  AN2 U3668 ( .A(n3521), .B(n3522), .Z(n3517) );
  AN2 U3669 ( .A(N4851), .B(N4831), .Z(n3522) );
  AN2 U3670 ( .A(N4941), .B(N4921), .Z(n3521) );
  AN2 U3671 ( .A(n3523), .B(n3524), .Z(n3507) );
  AN2 U3672 ( .A(n3525), .B(n3526), .Z(n3524) );
  AN2 U3673 ( .A(n3527), .B(n3528), .Z(n3526) );
  AN2 U3674 ( .A(N4981), .B(N4961), .Z(n3528) );
  AN2 U3675 ( .A(N5021), .B(N5001), .Z(n3527) );
  AN2 U3676 ( .A(n3529), .B(n3530), .Z(n3525) );
  AN2 U3677 ( .A(N5122), .B(N5102), .Z(n3530) );
  AN2 U3678 ( .A(N5251), .B(N5161), .Z(n3529) );
  AN2 U3679 ( .A(n3531), .B(n3532), .Z(n3523) );
  AN2 U3680 ( .A(n3533), .B(n3534), .Z(n3532) );
  AN2 U3681 ( .A(N5291), .B(N5271), .Z(n3534) );
  AN2 U3682 ( .A(N5610), .B(N5341), .Z(n3533) );
  AN2 U3683 ( .A(n3535), .B(N9910), .Z(n3531) );
  AN2 U3684 ( .A(N8010), .B(N7810), .Z(n3535) );
  IV U3685 ( .A(n3536), .Z(n147) );
  AN2 U3686 ( .A(n3537), .B(n3538), .Z(n3536) );
  AN2 U3687 ( .A(n3539), .B(n3540), .Z(n3538) );
  AN2 U3688 ( .A(n3541), .B(n3542), .Z(n3540) );
  AN2 U3689 ( .A(n3543), .B(n3544), .Z(n3542) );
  AN2 U3690 ( .A(n3545), .B(n3546), .Z(n3544) );
  AN2 U3691 ( .A(n3547), .B(n3548), .Z(n3546) );
  AN2 U3692 ( .A(N10310), .B(n3549), .Z(n3548) );
  IV U3693 ( .A(N6971), .Z(n3549) );
  AN2 U3694 ( .A(N10910), .B(N10510), .Z(n3547) );
  AN2 U3695 ( .A(n3550), .B(n3551), .Z(n3545) );
  AN2 U3696 ( .A(N1212), .B(N1192), .Z(n3551) );
  AN2 U3697 ( .A(N1271), .B(N1231), .Z(n3550) );
  AN2 U3698 ( .A(n3552), .B(n3553), .Z(n3543) );
  AN2 U3699 ( .A(n3554), .B(n3555), .Z(n3553) );
  AN2 U3700 ( .A(N1512), .B(N1361), .Z(n3555) );
  AN2 U3701 ( .A(N1691), .B(N1551), .Z(n3554) );
  AN2 U3702 ( .A(n3556), .B(n3557), .Z(n3552) );
  AN2 U3703 ( .A(N1771), .B(N1712), .Z(n3557) );
  AN2 U3704 ( .A(N1831), .B(N1812), .Z(n3556) );
  AN2 U3705 ( .A(n3558), .B(n3559), .Z(n3541) );
  AN2 U3706 ( .A(n3560), .B(n3561), .Z(n3559) );
  AN2 U3707 ( .A(n3562), .B(n3563), .Z(n3561) );
  AN2 U3708 ( .A(N1891), .B(N1851), .Z(n3563) );
  AN2 U3709 ( .A(N1931), .B(N1912), .Z(n3562) );
  AN2 U3710 ( .A(n3564), .B(n3565), .Z(n3560) );
  AN2 U3711 ( .A(N2051), .B(N1971), .Z(n3565) );
  AN2 U3712 ( .A(N2221), .B(N2191), .Z(n3564) );
  AN2 U3713 ( .A(n3566), .B(n3567), .Z(n3558) );
  AN2 U3714 ( .A(n3568), .B(n3569), .Z(n3567) );
  AN2 U3715 ( .A(N2381), .B(N2361), .Z(n3569) );
  AN2 U3716 ( .A(N2481), .B(N2441), .Z(n3568) );
  AN2 U3717 ( .A(n3570), .B(N2551), .Z(n3566) );
  AN2 U3718 ( .A(N2521), .B(N2501), .Z(n3570) );
  AN2 U3719 ( .A(n3571), .B(n3572), .Z(n3539) );
  AN2 U3720 ( .A(n3573), .B(n3574), .Z(n3572) );
  AN2 U3721 ( .A(n3575), .B(n3576), .Z(n3574) );
  AN2 U3722 ( .A(n3577), .B(n3578), .Z(n3576) );
  AN2 U3723 ( .A(N2591), .B(N2571), .Z(n3578) );
  AN2 U3724 ( .A(N2712), .B(N2631), .Z(n3577) );
  AN2 U3725 ( .A(n3579), .B(n3580), .Z(n3575) );
  AN2 U3726 ( .A(N2881), .B(N2851), .Z(n3580) );
  AN2 U3727 ( .A(N3041), .B(N3021), .Z(n3579) );
  AN2 U3728 ( .A(n3581), .B(n3582), .Z(n3573) );
  AN2 U3729 ( .A(n3583), .B(n3584), .Z(n3582) );
  AN2 U3730 ( .A(N3142), .B(N3102), .Z(n3584) );
  AN2 U3731 ( .A(N3181), .B(N3161), .Z(n3583) );
  AN2 U3732 ( .A(n3585), .B(N3341), .Z(n3581) );
  AN2 U3733 ( .A(N3321), .B(N3281), .Z(n3585) );
  AN2 U3734 ( .A(n3586), .B(n3587), .Z(n3571) );
  AN2 U3735 ( .A(n3588), .B(n3589), .Z(n3587) );
  AN2 U3736 ( .A(n3590), .B(n3591), .Z(n3589) );
  AN2 U3737 ( .A(N3401), .B(N3361), .Z(n3591) );
  AN2 U3738 ( .A(N3441), .B(N3421), .Z(n3590) );
  AN2 U3739 ( .A(n3592), .B(n3593), .Z(n3588) );
  AN2 U3740 ( .A(N3481), .B(N3461), .Z(n3593) );
  AN2 U3741 ( .A(N3571), .B(N3501), .Z(n3592) );
  AN2 U3742 ( .A(n3594), .B(n3595), .Z(n3586) );
  AN2 U3743 ( .A(n3596), .B(n3597), .Z(n3595) );
  AN2 U3744 ( .A(N3612), .B(N3591), .Z(n3597) );
  AN2 U3745 ( .A(N3651), .B(N3631), .Z(n3596) );
  AN2 U3746 ( .A(n3598), .B(N3751), .Z(n3594) );
  AN2 U3747 ( .A(N3731), .B(N3671), .Z(n3598) );
  AN2 U3748 ( .A(n3599), .B(n3600), .Z(n3537) );
  AN2 U3749 ( .A(n3601), .B(n3602), .Z(n3600) );
  AN2 U3750 ( .A(n3603), .B(n3604), .Z(n3602) );
  AN2 U3751 ( .A(n3605), .B(n3606), .Z(n3604) );
  AN2 U3752 ( .A(n3607), .B(n3608), .Z(n3606) );
  AN2 U3753 ( .A(N3881), .B(N3791), .Z(n3608) );
  AN2 U3754 ( .A(N3921), .B(N3901), .Z(n3607) );
  AN2 U3755 ( .A(n3609), .B(n3610), .Z(n3605) );
  AN2 U3756 ( .A(N4010), .B(N3961), .Z(n3610) );
  AN2 U3757 ( .A(N4181), .B(N4041), .Z(n3609) );
  AN2 U3758 ( .A(n3611), .B(n3612), .Z(n3603) );
  AN2 U3759 ( .A(n3613), .B(n3614), .Z(n3612) );
  AN2 U3760 ( .A(N4351), .B(N4212), .Z(n3614) );
  AN2 U3761 ( .A(N4431), .B(N4371), .Z(n3613) );
  AN2 U3762 ( .A(n3615), .B(N4512), .Z(n3611) );
  AN2 U3763 ( .A(N4491), .B(N4471), .Z(n3615) );
  AN2 U3764 ( .A(n3616), .B(n3617), .Z(n3601) );
  AN2 U3765 ( .A(n3618), .B(n3619), .Z(n3617) );
  AN2 U3766 ( .A(n3620), .B(n3621), .Z(n3619) );
  AN2 U3767 ( .A(N4571), .B(N4551), .Z(n3621) );
  AN2 U3768 ( .A(N4631), .B(N4591), .Z(n3620) );
  AN2 U3769 ( .A(n3622), .B(n3623), .Z(n3618) );
  AN2 U3770 ( .A(N4721), .B(N4710), .Z(n3623) );
  AN2 U3771 ( .A(N4901), .B(N4871), .Z(n3622) );
  AN2 U3772 ( .A(n3624), .B(n3625), .Z(n3616) );
  AN2 U3773 ( .A(n3626), .B(n3627), .Z(n3625) );
  AN2 U3774 ( .A(N5081), .B(N5061), .Z(n3627) );
  AN2 U3775 ( .A(N5141), .B(N5110), .Z(n3626) );
  AN2 U3776 ( .A(n3628), .B(N5221), .Z(n3624) );
  AN2 U3777 ( .A(N5201), .B(N5181), .Z(n3628) );
  AN2 U3778 ( .A(n3629), .B(n3630), .Z(n3599) );
  AN2 U3779 ( .A(n3631), .B(n3632), .Z(n3630) );
  AN2 U3780 ( .A(n3633), .B(n3634), .Z(n3632) );
  AN2 U3781 ( .A(n3635), .B(n3636), .Z(n3634) );
  AN2 U3782 ( .A(N5371), .B(N5321), .Z(n3636) );
  AN2 U3783 ( .A(N5410), .B(N5401), .Z(n3635) );
  AN2 U3784 ( .A(n3637), .B(n3638), .Z(n3633) );
  AN2 U3785 ( .A(N5531), .B(N5421), .Z(n3638) );
  AN2 U3786 ( .A(N5581), .B(N5561), .Z(n3637) );
  AN2 U3787 ( .A(n3639), .B(n3640), .Z(n3631) );
  AN2 U3788 ( .A(n3641), .B(n3642), .Z(n3640) );
  AN2 U3789 ( .A(N5631), .B(N5612), .Z(n3642) );
  AN2 U3790 ( .A(N5791), .B(N5651), .Z(n3641) );
  AN2 U3791 ( .A(n3643), .B(N5871), .Z(n3639) );
  AN2 U3792 ( .A(N5841), .B(N5821), .Z(n3643) );
  AN2 U3793 ( .A(n3644), .B(n3645), .Z(n3629) );
  AN2 U3794 ( .A(n3646), .B(n3647), .Z(n3645) );
  AN2 U3795 ( .A(n3648), .B(n3649), .Z(n3647) );
  AN2 U3796 ( .A(N5912), .B(N5891), .Z(n3649) );
  AN2 U3797 ( .A(N6010), .B(N5991), .Z(n3648) );
  AN2 U3798 ( .A(n3650), .B(n3651), .Z(n3646) );
  AN2 U3799 ( .A(N6610), .B(N6310), .Z(n3651) );
  AN2 U3800 ( .A(N7310), .B(N7010), .Z(n3650) );
  AN2 U3801 ( .A(n3652), .B(n3653), .Z(n3644) );
  AN2 U3802 ( .A(n3654), .B(n3655), .Z(n3653) );
  AN2 U3803 ( .A(N8510), .B(N7610), .Z(n3655) );
  AN2 U3804 ( .A(N9010), .B(N8810), .Z(n3654) );
  AN2 U3805 ( .A(n3656), .B(N9710), .Z(n3652) );
  AN2 U3806 ( .A(N9510), .B(N9310), .Z(n3656) );
  IV U3807 ( .A(N246), .Z(n145) );
  IV U3808 ( .A(N10), .Z(n14) );
  IV U3809 ( .A(N468), .Z(n139) );
  IV U3810 ( .A(N536), .Z(n137) );
  IV U3811 ( .A(tx_enc_sel[0]), .Z(n13) );
  IV U3812 ( .A(tx_enc_sel[1]), .Z(n12) );
  IV U3813 ( .A(tx_enc_sel[2]), .Z(n11) );
  IV U3814 ( .A(N324), .Z(n107) );
  IV U3815 ( .A(N526), .Z(n101) );
  IV U3816 ( .A(N86), .Z(n10) );
  IV U3817 ( .A(N91), .Z(n1) );
  OR2 U3818 ( .A(n3657), .B(n3658), .Z(N976) );
  OR2 U3819 ( .A(n3659), .B(n3660), .Z(n3658) );
  OR2 U3820 ( .A(n3661), .B(n3662), .Z(n3660) );
  OR2 U3821 ( .A(n3663), .B(n3664), .Z(n3657) );
  OR2 U3822 ( .A(N904), .B(n3665), .Z(n3663) );
  OR2 U3823 ( .A(n3666), .B(n3667), .Z(N955) );
  OR2 U3824 ( .A(n3668), .B(n3669), .Z(n3667) );
  OR2 U3825 ( .A(N922), .B(n20), .Z(n3666) );
  OR2 U3826 ( .A(n3670), .B(n3671), .Z(N952) );
  OR2 U3827 ( .A(n3668), .B(n3670), .Z(N932) );
  OR2 U3828 ( .A(n3672), .B(n3673), .Z(n3670) );
  OR2 U3829 ( .A(n3674), .B(n3675), .Z(n3673) );
  OR2 U3830 ( .A(n3676), .B(n3677), .Z(n3675) );
  OR2 U3831 ( .A(n3678), .B(n3679), .Z(n3677) );
  OR2 U3832 ( .A(n3680), .B(n3681), .Z(n3679) );
  OR2 U3833 ( .A(n3682), .B(n3683), .Z(n3678) );
  OR2 U3834 ( .A(n3684), .B(n3685), .Z(n3676) );
  OR2 U3835 ( .A(n3686), .B(n3687), .Z(n3685) );
  OR2 U3836 ( .A(n3688), .B(n3689), .Z(n3684) );
  OR2 U3837 ( .A(n3690), .B(n3691), .Z(n3674) );
  OR2 U3838 ( .A(n3692), .B(n3693), .Z(n3691) );
  OR2 U3839 ( .A(n3694), .B(n3695), .Z(n3693) );
  OR2 U3840 ( .A(n3696), .B(n3697), .Z(n3692) );
  OR2 U3841 ( .A(n3698), .B(n3699), .Z(n3690) );
  OR2 U3842 ( .A(n3700), .B(n3701), .Z(n3699) );
  OR2 U3843 ( .A(n3702), .B(n3703), .Z(n3698) );
  OR2 U3844 ( .A(n3704), .B(n3705), .Z(n3672) );
  OR2 U3845 ( .A(n3706), .B(n3707), .Z(n3705) );
  OR2 U3846 ( .A(n3708), .B(n3709), .Z(n3707) );
  OR2 U3847 ( .A(n3710), .B(n3711), .Z(n3709) );
  OR2 U3848 ( .A(n155), .B(n133), .Z(n3708) );
  IV U3849 ( .A(N668), .Z(n133) );
  IV U3850 ( .A(N7311), .Z(n155) );
  OR2 U3851 ( .A(n3712), .B(n3713), .Z(n3706) );
  OR2 U3852 ( .A(n180), .B(n174), .Z(n3713) );
  IV U3853 ( .A(N719), .Z(n174) );
  IV U3854 ( .A(N7011), .Z(n180) );
  OR2 U3855 ( .A(n205), .B(n181), .Z(n3712) );
  IV U3856 ( .A(N666), .Z(n181) );
  IV U3857 ( .A(N683), .Z(n205) );
  OR2 U3858 ( .A(n3714), .B(n3715), .Z(n3704) );
  OR2 U3859 ( .A(n3716), .B(n3717), .Z(n3715) );
  OR2 U3860 ( .A(n218), .B(n21), .Z(n3717) );
  IV U3861 ( .A(N725), .Z(n21) );
  IV U3862 ( .A(N674), .Z(n218) );
  OR2 U3863 ( .A(n25), .B(n24), .Z(n3716) );
  IV U3864 ( .A(N733), .Z(n24) );
  IV U3865 ( .A(N698), .Z(n25) );
  OR2 U3866 ( .A(n3718), .B(n3719), .Z(n3714) );
  OR2 U3867 ( .A(n28), .B(n267), .Z(n3719) );
  IV U3868 ( .A(N670), .Z(n267) );
  IV U3869 ( .A(N717), .Z(n28) );
  OR2 U3870 ( .A(n35), .B(n29), .Z(n3718) );
  IV U3871 ( .A(N6811), .Z(n29) );
  IV U3872 ( .A(N729), .Z(n35) );
  OR2 U3873 ( .A(n3720), .B(n3721), .Z(n3668) );
  OR2 U3874 ( .A(n3722), .B(n3723), .Z(n3721) );
  OR2 U3875 ( .A(n3724), .B(n3725), .Z(n3723) );
  OR2 U3876 ( .A(n3726), .B(n3727), .Z(n3725) );
  OR2 U3877 ( .A(n3728), .B(n3729), .Z(n3727) );
  OR2 U3878 ( .A(n3730), .B(n3731), .Z(n3726) );
  OR2 U3879 ( .A(n3732), .B(n3733), .Z(n3724) );
  OR2 U3880 ( .A(n3734), .B(n3735), .Z(n3733) );
  OR2 U3881 ( .A(n3736), .B(n3737), .Z(n3732) );
  OR2 U3882 ( .A(n3738), .B(n3739), .Z(n3722) );
  OR2 U3883 ( .A(n3740), .B(n3741), .Z(n3739) );
  OR2 U3884 ( .A(n3742), .B(n3743), .Z(n3741) );
  OR2 U3885 ( .A(n3744), .B(n3745), .Z(n3740) );
  OR2 U3886 ( .A(n3746), .B(n3747), .Z(n3738) );
  OR2 U3887 ( .A(n3748), .B(n3749), .Z(n3747) );
  OR2 U3888 ( .A(n3750), .B(n3751), .Z(n3746) );
  OR2 U3889 ( .A(n3752), .B(n3753), .Z(n3720) );
  OR2 U3890 ( .A(n3754), .B(n3755), .Z(n3753) );
  OR2 U3891 ( .A(n3756), .B(n3757), .Z(n3755) );
  OR2 U3892 ( .A(n3758), .B(n3759), .Z(n3757) );
  OR2 U3893 ( .A(n182), .B(n135), .Z(n3756) );
  IV U3894 ( .A(N602), .Z(n135) );
  IV U3895 ( .A(N633), .Z(n182) );
  OR2 U3896 ( .A(n3760), .B(n3761), .Z(n3754) );
  OR2 U3897 ( .A(n206), .B(n183), .Z(n3761) );
  IV U3898 ( .A(N600), .Z(n183) );
  IV U3899 ( .A(N649), .Z(n206) );
  OR2 U3900 ( .A(n220), .B(n207), .Z(n3760) );
  IV U3901 ( .A(N616), .Z(n207) );
  IV U3902 ( .A(N608), .Z(n220) );
  OR2 U3903 ( .A(n3762), .B(n3763), .Z(n3752) );
  OR2 U3904 ( .A(n3764), .B(n3765), .Z(n3763) );
  OR2 U3905 ( .A(n269), .B(n231), .Z(n3765) );
  IV U3906 ( .A(N6611), .Z(n231) );
  IV U3907 ( .A(N604), .Z(n269) );
  OR2 U3908 ( .A(n60), .B(n48), .Z(n3764) );
  IV U3909 ( .A(N655), .Z(n48) );
  IV U3910 ( .A(N663), .Z(n60) );
  OR2 U3911 ( .A(n3766), .B(n3767), .Z(n3762) );
  OR2 U3912 ( .A(n72), .B(n61), .Z(n3767) );
  IV U3913 ( .A(N630), .Z(n61) );
  IV U3914 ( .A(N647), .Z(n72) );
  OR2 U3915 ( .A(n97), .B(n73), .Z(n3766) );
  IV U3916 ( .A(N614), .Z(n73) );
  IV U3917 ( .A(N659), .Z(n97) );
  OR2 U3918 ( .A(n3768), .B(n3769), .Z(N908) );
  OR2 U3919 ( .A(n3669), .B(n3671), .Z(n3769) );
  OR2 U3920 ( .A(n3770), .B(n3771), .Z(n3671) );
  OR2 U3921 ( .A(n3772), .B(n3773), .Z(n3771) );
  OR2 U3922 ( .A(n3774), .B(n3775), .Z(n3773) );
  OR2 U3923 ( .A(n3776), .B(n3777), .Z(n3775) );
  OR2 U3924 ( .A(n3778), .B(n3779), .Z(n3777) );
  OR2 U3925 ( .A(n3780), .B(n3781), .Z(n3776) );
  OR2 U3926 ( .A(n3782), .B(n3783), .Z(n3774) );
  OR2 U3927 ( .A(n3784), .B(n3785), .Z(n3783) );
  OR2 U3928 ( .A(n3786), .B(n3787), .Z(n3782) );
  OR2 U3929 ( .A(n3788), .B(n3789), .Z(n3772) );
  OR2 U3930 ( .A(n3790), .B(n3791), .Z(n3789) );
  OR2 U3931 ( .A(n3792), .B(n3793), .Z(n3791) );
  OR2 U3932 ( .A(n3794), .B(n3795), .Z(n3790) );
  OR2 U3933 ( .A(n3796), .B(n3797), .Z(n3788) );
  OR2 U3934 ( .A(n3798), .B(n3799), .Z(n3797) );
  OR2 U3935 ( .A(n3800), .B(n3801), .Z(n3796) );
  OR2 U3936 ( .A(n3802), .B(n3803), .Z(n3770) );
  OR2 U3937 ( .A(n3804), .B(n3805), .Z(n3803) );
  OR2 U3938 ( .A(n3806), .B(n3807), .Z(n3805) );
  OR2 U3939 ( .A(n3808), .B(n3809), .Z(n3807) );
  OR2 U3940 ( .A(n141), .B(n103), .Z(n3806) );
  IV U3941 ( .A(N457), .Z(n103) );
  IV U3942 ( .A(N400), .Z(n141) );
  OR2 U3943 ( .A(n3810), .B(n3811), .Z(n3804) );
  OR2 U3944 ( .A(n189), .B(n188), .Z(n3811) );
  IV U3945 ( .A(N4311), .Z(n188) );
  IV U3946 ( .A(N398), .Z(n189) );
  OR2 U3947 ( .A(n213), .B(n212), .Z(n3810) );
  IV U3948 ( .A(N447), .Z(n212) );
  IV U3949 ( .A(N414), .Z(n213) );
  OR2 U3950 ( .A(n3812), .B(n3813), .Z(n3802) );
  OR2 U3951 ( .A(n3814), .B(n3815), .Z(n3813) );
  OR2 U3952 ( .A(n237), .B(n226), .Z(n3815) );
  IV U3953 ( .A(N406), .Z(n226) );
  IV U3954 ( .A(N459), .Z(n237) );
  OR2 U3955 ( .A(n54), .B(n275), .Z(n3814) );
  IV U3956 ( .A(N402), .Z(n275) );
  IV U3957 ( .A(N453), .Z(n54) );
  OR2 U3958 ( .A(n3816), .B(n3817), .Z(n3812) );
  OR2 U3959 ( .A(n67), .B(n66), .Z(n3817) );
  IV U3960 ( .A(N4611), .Z(n66) );
  IV U3961 ( .A(N428), .Z(n67) );
  OR2 U3962 ( .A(n79), .B(n78), .Z(n3816) );
  IV U3963 ( .A(N445), .Z(n78) );
  IV U3964 ( .A(N4121), .Z(n79) );
  OR2 U3965 ( .A(n3818), .B(n3819), .Z(n3669) );
  OR2 U3966 ( .A(n3820), .B(n3821), .Z(n3819) );
  OR2 U3967 ( .A(n3822), .B(n3823), .Z(n3821) );
  OR2 U3968 ( .A(n3824), .B(n3825), .Z(n3823) );
  OR2 U3969 ( .A(n3826), .B(n3827), .Z(n3825) );
  OR2 U3970 ( .A(n3828), .B(n3829), .Z(n3824) );
  OR2 U3971 ( .A(n3830), .B(n3831), .Z(n3822) );
  OR2 U3972 ( .A(n3832), .B(n3833), .Z(n3831) );
  OR2 U3973 ( .A(n3834), .B(n3835), .Z(n3830) );
  OR2 U3974 ( .A(n3836), .B(n3837), .Z(n3820) );
  OR2 U3975 ( .A(n3838), .B(n3839), .Z(n3837) );
  OR2 U3976 ( .A(n3840), .B(n3841), .Z(n3839) );
  OR2 U3977 ( .A(n3842), .B(n3843), .Z(n3838) );
  OR2 U3978 ( .A(n3844), .B(n3845), .Z(n3836) );
  OR2 U3979 ( .A(n3846), .B(n3847), .Z(n3845) );
  OR2 U3980 ( .A(n3848), .B(n3849), .Z(n3844) );
  OR2 U3981 ( .A(n3850), .B(n3851), .Z(n3818) );
  OR2 U3982 ( .A(n3852), .B(n3853), .Z(n3851) );
  OR2 U3983 ( .A(n3854), .B(n3855), .Z(n3853) );
  OR2 U3984 ( .A(n3856), .B(n3857), .Z(n3855) );
  OR2 U3985 ( .A(n143), .B(n105), .Z(n3854) );
  IV U3986 ( .A(N3911), .Z(n105) );
  IV U3987 ( .A(N334), .Z(n143) );
  OR2 U3988 ( .A(n3858), .B(n3859), .Z(n3852) );
  OR2 U3989 ( .A(n191), .B(n190), .Z(n3859) );
  IV U3990 ( .A(N365), .Z(n190) );
  IV U3991 ( .A(N332), .Z(n191) );
  OR2 U3992 ( .A(n215), .B(n214), .Z(n3858) );
  IV U3993 ( .A(N3811), .Z(n214) );
  IV U3994 ( .A(N348), .Z(n215) );
  OR2 U3995 ( .A(n3860), .B(n3861), .Z(n3850) );
  OR2 U3996 ( .A(n3862), .B(n3863), .Z(n3861) );
  OR2 U3997 ( .A(n239), .B(n228), .Z(n3863) );
  IV U3998 ( .A(N340), .Z(n228) );
  IV U3999 ( .A(N393), .Z(n239) );
  OR2 U4000 ( .A(n56), .B(n277), .Z(n3862) );
  IV U4001 ( .A(N336), .Z(n277) );
  IV U4002 ( .A(N387), .Z(n56) );
  OR2 U4003 ( .A(n3864), .B(n3865), .Z(n3860) );
  OR2 U4004 ( .A(n69), .B(n68), .Z(n3865) );
  IV U4005 ( .A(N395), .Z(n68) );
  IV U4006 ( .A(N362), .Z(n69) );
  OR2 U4007 ( .A(n81), .B(n80), .Z(n3864) );
  IV U4008 ( .A(N379), .Z(n80) );
  IV U4009 ( .A(N346), .Z(n81) );
  OR2 U4010 ( .A(N904), .B(n43), .Z(n3768) );
  OR2 U4011 ( .A(n3866), .B(n3867), .Z(N6641) );
  IV U4012 ( .A(n3868), .Z(n3867) );
  AN2 U4013 ( .A(N6141), .B(N6102), .Z(n3868) );
  OR2 U4014 ( .A(N6221), .B(n3869), .Z(n3866) );
  IV U4015 ( .A(N6041), .Z(n3869) );
  OR2 U4016 ( .A(n3870), .B(n3871), .Z(N6361) );
  OR2 U4017 ( .A(N6271), .B(N6261), .Z(n3871) );
  OR2 U4018 ( .A(N6281), .B(n3872), .Z(n3870) );
  OR2 U4019 ( .A(N6301), .B(N6291), .Z(n3872) );
  OR2 U4020 ( .A(N6241), .B(n3873), .Z(N6351) );
  OR2 U4021 ( .A(N6321), .B(N6251), .Z(n3873) );
  OR2 U4022 ( .A(n292), .B(n3874), .Z(N11811) );
  OR2 U4023 ( .A(n299), .B(n294), .Z(n3874) );
  IV U4024 ( .A(N845), .Z(n294) );
  IV U4025 ( .A(N855), .Z(n299) );
  IV U4026 ( .A(N870), .Z(n292) );
  OR2 U4027 ( .A(n3875), .B(n3876), .Z(N1158) );
  OR2 U4028 ( .A(n3877), .B(n3878), .Z(n3876) );
  OR2 U4029 ( .A(n3879), .B(n3880), .Z(n3878) );
  OR2 U4030 ( .A(n3881), .B(n3882), .Z(n3875) );
  OR2 U4031 ( .A(n3883), .B(n3884), .Z(n3882) );
  OR2 U4032 ( .A(N1154), .B(n3665), .Z(n3881) );
  OR2 U4033 ( .A(n3885), .B(n3886), .Z(n3665) );
  OR2 U4034 ( .A(n3887), .B(n3888), .Z(n3886) );
  OR2 U4035 ( .A(n3889), .B(n3890), .Z(n3885) );
  OR2 U4036 ( .A(n3891), .B(n3892), .Z(N1120) );
  OR2 U4037 ( .A(n3893), .B(n3894), .Z(n3892) );
  OR2 U4038 ( .A(n3895), .B(n3896), .Z(n3894) );
  OR2 U4039 ( .A(n3897), .B(n3898), .Z(n3891) );
  OR2 U4040 ( .A(N1116), .B(n3889), .Z(n3898) );
  OR2 U4041 ( .A(n3899), .B(n3900), .Z(n3889) );
  OR2 U4042 ( .A(n3901), .B(n3902), .Z(n3900) );
  OR2 U4043 ( .A(n3742), .B(n3694), .Z(n3902) );
  IV U4044 ( .A(N672), .Z(n3694) );
  IV U4045 ( .A(N606), .Z(n3742) );
  OR2 U4046 ( .A(n3840), .B(n3792), .Z(n3901) );
  IV U4047 ( .A(N404), .Z(n3792) );
  IV U4048 ( .A(N338), .Z(n3840) );
  OR2 U4049 ( .A(n3903), .B(n3904), .Z(n3899) );
  OR2 U4050 ( .A(n88), .B(n31), .Z(n3904) );
  IV U4051 ( .A(N7511), .Z(n31) );
  IV U4052 ( .A(N540), .Z(n88) );
  OR2 U4053 ( .A(n96), .B(n90), .Z(n3903) );
  IV U4054 ( .A(N472), .Z(n90) );
  IV U4055 ( .A(N253), .Z(n96) );
  OR2 U4056 ( .A(n3905), .B(n3906), .Z(N11011) );
  OR2 U4057 ( .A(n3907), .B(n3908), .Z(n3906) );
  OR2 U4058 ( .A(n3884), .B(n3909), .Z(n3908) );
  OR2 U4059 ( .A(n3910), .B(n3664), .Z(n3905) );
  OR2 U4060 ( .A(n3897), .B(n3911), .Z(n3664) );
  OR2 U4061 ( .A(n3912), .B(n3913), .Z(n3897) );
  OR2 U4062 ( .A(n3914), .B(n3915), .Z(n3913) );
  OR2 U4063 ( .A(n3748), .B(n3700), .Z(n3915) );
  IV U4064 ( .A(N679), .Z(n3700) );
  IV U4065 ( .A(N6121), .Z(n3748) );
  OR2 U4066 ( .A(n3846), .B(n3798), .Z(n3914) );
  IV U4067 ( .A(N4101), .Z(n3798) );
  IV U4068 ( .A(N344), .Z(n3846) );
  OR2 U4069 ( .A(n3916), .B(n3917), .Z(n3912) );
  OR2 U4070 ( .A(n258), .B(n162), .Z(n3917) );
  IV U4071 ( .A(N7611), .Z(n162) );
  IV U4072 ( .A(N546), .Z(n258) );
  OR2 U4073 ( .A(n266), .B(n260), .Z(n3916) );
  IV U4074 ( .A(N478), .Z(n260) );
  IV U4075 ( .A(N264), .Z(n266) );
  OR2 U4076 ( .A(N1097), .B(n3890), .Z(n3910) );
  OR2 U4077 ( .A(n3918), .B(n3919), .Z(n3890) );
  OR2 U4078 ( .A(n3920), .B(n3921), .Z(n3919) );
  OR2 U4079 ( .A(n3745), .B(n3697), .Z(n3921) );
  IV U4080 ( .A(N677), .Z(n3697) );
  IV U4081 ( .A(N6101), .Z(n3745) );
  OR2 U4082 ( .A(n3843), .B(n3795), .Z(n3920) );
  IV U4083 ( .A(N408), .Z(n3795) );
  IV U4084 ( .A(N342), .Z(n3843) );
  OR2 U4085 ( .A(n3922), .B(n3923), .Z(n3918) );
  OR2 U4086 ( .A(n126), .B(n124), .Z(n3923) );
  IV U4087 ( .A(N544), .Z(n124) );
  IV U4088 ( .A(N476), .Z(n126) );
  OR2 U4089 ( .A(n41), .B(n132), .Z(n3922) );
  IV U4090 ( .A(N2611), .Z(n132) );
  IV U4091 ( .A(N758), .Z(n41) );
  OR2 U4092 ( .A(n3924), .B(n3925), .Z(N1063) );
  OR2 U4093 ( .A(n3926), .B(n3927), .Z(n3925) );
  OR2 U4094 ( .A(n3895), .B(n3928), .Z(n3927) );
  OR2 U4095 ( .A(n3909), .B(n3929), .Z(n3895) );
  OR2 U4096 ( .A(n3661), .B(n3883), .Z(n3929) );
  OR2 U4097 ( .A(n3930), .B(n3931), .Z(n3883) );
  OR2 U4098 ( .A(n3932), .B(n3933), .Z(n3931) );
  OR2 U4099 ( .A(n3793), .B(n3695), .Z(n3933) );
  IV U4100 ( .A(N690), .Z(n3695) );
  IV U4101 ( .A(N420), .Z(n3793) );
  OR2 U4102 ( .A(n3841), .B(n3743), .Z(n3932) );
  IV U4103 ( .A(N622), .Z(n3743) );
  IV U4104 ( .A(N354), .Z(n3841) );
  OR2 U4105 ( .A(n3934), .B(n3935), .Z(n3930) );
  OR2 U4106 ( .A(n51), .B(n20), .Z(n3935) );
  IV U4107 ( .A(N777), .Z(n20) );
  IV U4108 ( .A(N556), .Z(n51) );
  OR2 U4109 ( .A(n59), .B(n53), .Z(n3934) );
  IV U4110 ( .A(N488), .Z(n53) );
  IV U4111 ( .A(N280), .Z(n59) );
  OR2 U4112 ( .A(n3936), .B(n3937), .Z(n3661) );
  OR2 U4113 ( .A(n3938), .B(n3939), .Z(n3937) );
  OR2 U4114 ( .A(n3750), .B(n3702), .Z(n3939) );
  IV U4115 ( .A(N688), .Z(n3702) );
  IV U4116 ( .A(N620), .Z(n3750) );
  OR2 U4117 ( .A(n3848), .B(n3800), .Z(n3938) );
  IV U4118 ( .A(N418), .Z(n3800) );
  IV U4119 ( .A(N352), .Z(n3848) );
  OR2 U4120 ( .A(n3940), .B(n3941), .Z(n3936) );
  OR2 U4121 ( .A(n246), .B(n158), .Z(n3941) );
  IV U4122 ( .A(N775), .Z(n158) );
  IV U4123 ( .A(N554), .Z(n246) );
  OR2 U4124 ( .A(n254), .B(n248), .Z(n3940) );
  IV U4125 ( .A(N486), .Z(n248) );
  IV U4126 ( .A(N278), .Z(n254) );
  OR2 U4127 ( .A(n3942), .B(n3943), .Z(n3909) );
  OR2 U4128 ( .A(n3944), .B(n3945), .Z(n3943) );
  OR2 U4129 ( .A(n3787), .B(n3689), .Z(n3945) );
  IV U4130 ( .A(N696), .Z(n3689) );
  IV U4131 ( .A(N426), .Z(n3787) );
  OR2 U4132 ( .A(n3835), .B(n3737), .Z(n3944) );
  IV U4133 ( .A(N628), .Z(n3737) );
  IV U4134 ( .A(N360), .Z(n3835) );
  OR2 U4135 ( .A(n3946), .B(n3947), .Z(n3942) );
  OR2 U4136 ( .A(n234), .B(n154), .Z(n3947) );
  IV U4137 ( .A(N784), .Z(n154) );
  IV U4138 ( .A(N562), .Z(n234) );
  OR2 U4139 ( .A(n242), .B(n236), .Z(n3946) );
  IV U4140 ( .A(N494), .Z(n236) );
  IV U4141 ( .A(N287), .Z(n242) );
  OR2 U4142 ( .A(n3948), .B(n3949), .Z(n3924) );
  OR2 U4143 ( .A(n3884), .B(n3950), .Z(n3949) );
  OR2 U4144 ( .A(n3951), .B(n3952), .Z(n3884) );
  OR2 U4145 ( .A(n3953), .B(n3954), .Z(n3952) );
  OR2 U4146 ( .A(n3786), .B(n3688), .Z(n3954) );
  IV U4147 ( .A(N694), .Z(n3688) );
  IV U4148 ( .A(N424), .Z(n3786) );
  OR2 U4149 ( .A(n3834), .B(n3736), .Z(n3953) );
  IV U4150 ( .A(N626), .Z(n3736) );
  IV U4151 ( .A(N358), .Z(n3834) );
  OR2 U4152 ( .A(n3955), .B(n3956), .Z(n3951) );
  OR2 U4153 ( .A(n102), .B(n100), .Z(n3956) );
  IV U4154 ( .A(N560), .Z(n100) );
  IV U4155 ( .A(N492), .Z(n102) );
  OR2 U4156 ( .A(n34), .B(n108), .Z(n3955) );
  IV U4157 ( .A(N285), .Z(n108) );
  IV U4158 ( .A(N782), .Z(n34) );
  OR2 U4159 ( .A(n3887), .B(n3911), .Z(n3948) );
  OR2 U4160 ( .A(n3957), .B(n3958), .Z(n3911) );
  OR2 U4161 ( .A(n3959), .B(n3960), .Z(n3958) );
  OR2 U4162 ( .A(n3751), .B(n3703), .Z(n3960) );
  IV U4163 ( .A(N692), .Z(n3703) );
  IV U4164 ( .A(N624), .Z(n3751) );
  OR2 U4165 ( .A(n3849), .B(n3801), .Z(n3959) );
  IV U4166 ( .A(N422), .Z(n3801) );
  IV U4167 ( .A(N356), .Z(n3849) );
  OR2 U4168 ( .A(n3961), .B(n3962), .Z(n3957) );
  OR2 U4169 ( .A(n196), .B(n169), .Z(n3962) );
  IV U4170 ( .A(N780), .Z(n169) );
  IV U4171 ( .A(N558), .Z(n196) );
  OR2 U4172 ( .A(n204), .B(n198), .Z(n3961) );
  IV U4173 ( .A(N490), .Z(n198) );
  IV U4174 ( .A(N283), .Z(n204) );
  OR2 U4175 ( .A(n3963), .B(n3964), .Z(n3887) );
  OR2 U4176 ( .A(n3965), .B(n3966), .Z(n3964) );
  OR2 U4177 ( .A(n3744), .B(n3696), .Z(n3966) );
  IV U4178 ( .A(N686), .Z(n3696) );
  IV U4179 ( .A(N618), .Z(n3744) );
  OR2 U4180 ( .A(n3842), .B(n3794), .Z(n3965) );
  IV U4181 ( .A(N416), .Z(n3794) );
  IV U4182 ( .A(N350), .Z(n3842) );
  OR2 U4183 ( .A(n3967), .B(n3968), .Z(n3963) );
  OR2 U4184 ( .A(n114), .B(n112), .Z(n3968) );
  IV U4185 ( .A(N552), .Z(n112) );
  IV U4186 ( .A(N484), .Z(n114) );
  OR2 U4187 ( .A(n38), .B(n120), .Z(n3967) );
  IV U4188 ( .A(N275), .Z(n120) );
  IV U4189 ( .A(N772), .Z(n38) );
  OR2 U4190 ( .A(n3969), .B(n3970), .Z(N1027) );
  OR2 U4191 ( .A(n3907), .B(n3926), .Z(n3970) );
  OR2 U4192 ( .A(n3877), .B(n3971), .Z(n3926) );
  OR2 U4193 ( .A(N9911), .B(n37), .Z(n3971) );
  IV U4194 ( .A(N8101), .Z(n37) );
  OR2 U4195 ( .A(n3972), .B(n3973), .Z(n3877) );
  OR2 U4196 ( .A(n3683), .B(n3974), .Z(n3973) );
  OR2 U4197 ( .A(n3731), .B(n3781), .Z(n3974) );
  IV U4198 ( .A(N449), .Z(n3781) );
  IV U4199 ( .A(N6511), .Z(n3731) );
  IV U4200 ( .A(N7211), .Z(n3683) );
  OR2 U4201 ( .A(n3975), .B(n3976), .Z(n3972) );
  OR2 U4202 ( .A(n111), .B(n3829), .Z(n3976) );
  IV U4203 ( .A(N383), .Z(n3829) );
  IV U4204 ( .A(N585), .Z(n111) );
  OR2 U4205 ( .A(n119), .B(n113), .Z(n3975) );
  IV U4206 ( .A(N518), .Z(n113) );
  IV U4207 ( .A(N3141), .Z(n119) );
  OR2 U4208 ( .A(n3977), .B(n3978), .Z(n3907) );
  OR2 U4209 ( .A(n3928), .B(n3979), .Z(n3978) );
  OR2 U4210 ( .A(n3879), .B(n3893), .Z(n3979) );
  OR2 U4211 ( .A(n3980), .B(n3981), .Z(n3893) );
  OR2 U4212 ( .A(n3682), .B(n3982), .Z(n3981) );
  OR2 U4213 ( .A(n3730), .B(n3780), .Z(n3982) );
  IV U4214 ( .A(N443), .Z(n3780) );
  IV U4215 ( .A(N645), .Z(n3730) );
  IV U4216 ( .A(N715), .Z(n3682) );
  OR2 U4217 ( .A(n3983), .B(n3984), .Z(n3980) );
  OR2 U4218 ( .A(n257), .B(n3828), .Z(n3984) );
  IV U4219 ( .A(N377), .Z(n3828) );
  IV U4220 ( .A(N579), .Z(n257) );
  OR2 U4221 ( .A(n265), .B(n259), .Z(n3983) );
  IV U4222 ( .A(N5121), .Z(n259) );
  IV U4223 ( .A(N308), .Z(n265) );
  OR2 U4224 ( .A(n3985), .B(n3986), .Z(n3879) );
  OR2 U4225 ( .A(n3687), .B(n3987), .Z(n3986) );
  OR2 U4226 ( .A(n3735), .B(n3785), .Z(n3987) );
  IV U4227 ( .A(N4411), .Z(n3785) );
  IV U4228 ( .A(N643), .Z(n3735) );
  IV U4229 ( .A(N7131), .Z(n3687) );
  OR2 U4230 ( .A(n3988), .B(n3989), .Z(n3985) );
  OR2 U4231 ( .A(n123), .B(n3833), .Z(n3989) );
  IV U4232 ( .A(N375), .Z(n3833) );
  IV U4233 ( .A(N577), .Z(n123) );
  OR2 U4234 ( .A(n131), .B(n125), .Z(n3988) );
  IV U4235 ( .A(N5101), .Z(n125) );
  IV U4236 ( .A(N306), .Z(n131) );
  OR2 U4237 ( .A(n3990), .B(n3991), .Z(n3928) );
  OR2 U4238 ( .A(n3681), .B(n3992), .Z(n3991) );
  OR2 U4239 ( .A(n3729), .B(n3779), .Z(n3992) );
  IV U4240 ( .A(N455), .Z(n3779) );
  IV U4241 ( .A(N657), .Z(n3729) );
  IV U4242 ( .A(N727), .Z(n3681) );
  OR2 U4243 ( .A(n3993), .B(n3994), .Z(n3990) );
  OR2 U4244 ( .A(n195), .B(n3827), .Z(n3994) );
  IV U4245 ( .A(N389), .Z(n3827) );
  IV U4246 ( .A(N5911), .Z(n195) );
  OR2 U4247 ( .A(n203), .B(n197), .Z(n3993) );
  IV U4248 ( .A(N524), .Z(n197) );
  IV U4249 ( .A(N3211), .Z(n203) );
  OR2 U4250 ( .A(n3662), .B(n3995), .Z(n3977) );
  OR2 U4251 ( .A(n40), .B(n175), .Z(n3995) );
  IV U4252 ( .A(N800), .Z(n175) );
  IV U4253 ( .A(N802), .Z(n40) );
  OR2 U4254 ( .A(n3996), .B(n3997), .Z(n3662) );
  OR2 U4255 ( .A(n3711), .B(n3998), .Z(n3997) );
  OR2 U4256 ( .A(n3809), .B(n3759), .Z(n3998) );
  IV U4257 ( .A(N6411), .Z(n3759) );
  IV U4258 ( .A(N439), .Z(n3809) );
  IV U4259 ( .A(N7111), .Z(n3711) );
  OR2 U4260 ( .A(n3999), .B(n4000), .Z(n3996) );
  OR2 U4261 ( .A(n221), .B(n3857), .Z(n4000) );
  IV U4262 ( .A(N373), .Z(n3857) );
  IV U4263 ( .A(N575), .Z(n221) );
  OR2 U4264 ( .A(n229), .B(n223), .Z(n3999) );
  IV U4265 ( .A(N508), .Z(n223) );
  IV U4266 ( .A(N304), .Z(n229) );
  OR2 U4267 ( .A(n3896), .B(n4001), .Z(n3969) );
  OR2 U4268 ( .A(n161), .B(n3888), .Z(n4001) );
  OR2 U4269 ( .A(n4002), .B(n4003), .Z(n3888) );
  OR2 U4270 ( .A(n4004), .B(n4005), .Z(n4003) );
  OR2 U4271 ( .A(n3749), .B(n3701), .Z(n4005) );
  IV U4272 ( .A(N703), .Z(n3701) );
  IV U4273 ( .A(N635), .Z(n3749) );
  OR2 U4274 ( .A(n3847), .B(n3799), .Z(n4004) );
  IV U4275 ( .A(N433), .Z(n3799) );
  IV U4276 ( .A(N367), .Z(n3847) );
  OR2 U4277 ( .A(n4006), .B(n4007), .Z(n4002) );
  OR2 U4278 ( .A(n138), .B(n136), .Z(n4007) );
  IV U4279 ( .A(N569), .Z(n136) );
  IV U4280 ( .A(N502), .Z(n138) );
  OR2 U4281 ( .A(n43), .B(n144), .Z(n4006) );
  IV U4282 ( .A(N298), .Z(n144) );
  IV U4283 ( .A(N794), .Z(n43) );
  IV U4284 ( .A(N804), .Z(n161) );
  OR2 U4285 ( .A(n4008), .B(n4009), .Z(n3896) );
  OR2 U4286 ( .A(n3880), .B(n3950), .Z(n4009) );
  OR2 U4287 ( .A(n4010), .B(n4011), .Z(n3950) );
  OR2 U4288 ( .A(n3680), .B(n4012), .Z(n4011) );
  OR2 U4289 ( .A(n3728), .B(n3778), .Z(n4012) );
  IV U4290 ( .A(N4511), .Z(n3778) );
  IV U4291 ( .A(N653), .Z(n3728) );
  IV U4292 ( .A(N723), .Z(n3680) );
  OR2 U4293 ( .A(n4013), .B(n4014), .Z(n4010) );
  OR2 U4294 ( .A(n245), .B(n3826), .Z(n4014) );
  IV U4295 ( .A(N385), .Z(n3826) );
  IV U4296 ( .A(N587), .Z(n245) );
  OR2 U4297 ( .A(n253), .B(n247), .Z(n4013) );
  IV U4298 ( .A(N520), .Z(n247) );
  IV U4299 ( .A(N316), .Z(n253) );
  OR2 U4300 ( .A(n4015), .B(n4016), .Z(n3880) );
  OR2 U4301 ( .A(n4017), .B(n4018), .Z(n4016) );
  OR2 U4302 ( .A(n3784), .B(n3686), .Z(n4018) );
  IV U4303 ( .A(N709), .Z(n3686) );
  IV U4304 ( .A(N437), .Z(n3784) );
  OR2 U4305 ( .A(n3832), .B(n3734), .Z(n4017) );
  IV U4306 ( .A(N639), .Z(n3734) );
  IV U4307 ( .A(N3711), .Z(n3832) );
  OR2 U4308 ( .A(n4019), .B(n4020), .Z(n4015) );
  OR2 U4309 ( .A(n87), .B(n30), .Z(n4020) );
  IV U4310 ( .A(N798), .Z(n30) );
  IV U4311 ( .A(N573), .Z(n87) );
  OR2 U4312 ( .A(n95), .B(n89), .Z(n4019) );
  IV U4313 ( .A(N506), .Z(n89) );
  IV U4314 ( .A(N302), .Z(n95) );
  OR2 U4315 ( .A(n165), .B(n3659), .Z(n4008) );
  OR2 U4316 ( .A(n4021), .B(n4022), .Z(n3659) );
  OR2 U4317 ( .A(n3710), .B(n4023), .Z(n4022) );
  OR2 U4318 ( .A(n3808), .B(n3758), .Z(n4023) );
  IV U4319 ( .A(N637), .Z(n3758) );
  IV U4320 ( .A(N435), .Z(n3808) );
  IV U4321 ( .A(N707), .Z(n3710) );
  OR2 U4322 ( .A(n4024), .B(n4025), .Z(n4021) );
  OR2 U4323 ( .A(n270), .B(n3856), .Z(n4025) );
  IV U4324 ( .A(N369), .Z(n3856) );
  IV U4325 ( .A(N5711), .Z(n270) );
  OR2 U4326 ( .A(n278), .B(n272), .Z(n4024) );
  IV U4327 ( .A(N504), .Z(n272) );
  IV U4328 ( .A(N300), .Z(n278) );
  IV U4329 ( .A(N796), .Z(n165) );
endmodule

