
module PCIEXP_TX ( PCLK250, RST_BeaconEnable_R0, CNTL_RESETN_P0, 
        CNTL_Loopback_P0, CNTL_TXEnable_P0, RX_LoopbackData_P2, TXCOMPLIANCE, 
        TXDATA, TXDATAK, TXELECIDLE, HSS_TXBEACONCMD, HSS_TXD, HSS_TXELECIDLE, 
        assertion_shengyushen );
  input [9:0] RX_LoopbackData_P2;
  input [7:0] TXDATA;
  output [9:0] HSS_TXD;
  input PCLK250, RST_BeaconEnable_R0, CNTL_RESETN_P0, CNTL_Loopback_P0,
         CNTL_TXEnable_P0, TXCOMPLIANCE, TXDATAK, TXELECIDLE;
  output HSS_TXBEACONCMD, HSS_TXELECIDLE, assertion_shengyushen;
  wire   n3, n4, n10, n11, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n25, n26, n28, n29, n30, n31, n32, n33, n35, n36, n37, n39, n40, n41,
         n44, n46, n48, n49, n52, n55, n58, n59, n60, n63, n64, n65, n68, n69,
         n71, n72, n73, n74, n76, n78, n80, n82, n84, n86, n87, n89, n91, n93,
         n94, n96, n97, n98, n100, n101, n102, n104, n105, n106, n108, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n140, n141, n142, n145, n146, n147,
         n148, n149, n150, n151, n153, n154, n157, n158, n159, n160, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n206, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, U6_Z_0,
         U6_DATA2_0, U5_DATA2_4, U5_DATA2_5, U4_Z_0, n351, n353, n354, n356,
         n358, n360, n362, n364, n366, n368, n370, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566;
  wire   [5:9] n;

  OR2 C36 ( .A(n426), .B(n427), .Z(n25) );
  OR2 C37 ( .A(n229), .B(n25), .Z(n26) );
  AN2 C39 ( .A(n223), .B(n222), .Z(n28) );
  AN2 C40 ( .A(n224), .B(n28), .Z(n29) );
  AN2 C41 ( .A(n225), .B(n29), .Z(n30) );
  OR2 C42 ( .A(n223), .B(n222), .Z(n31) );
  OR2 C43 ( .A(n224), .B(n31), .Z(n32) );
  OR2 C44 ( .A(n225), .B(n32), .Z(n33) );
  AN2 C46 ( .A(n228), .B(n227), .Z(n35) );
  AN2 C47 ( .A(n229), .B(n35), .Z(n36) );
  OR2 C48 ( .A(U5_DATA2_5), .B(U5_DATA2_4), .Z(n37) );
  AN2 C50 ( .A(U5_DATA2_5), .B(U5_DATA2_4), .Z(n39) );
  OR2 C53 ( .A(n228), .B(n227), .Z(n40) );
  OR2 C54 ( .A(n229), .B(n40), .Z(n41) );
  OR2 C58 ( .A(n423), .B(n40), .Z(n44) );
  OR2 C60 ( .A(n225), .B(n224), .Z(n46) );
  OR2 C67 ( .A(n446), .B(n68), .Z(n48) );
  OR2 C68 ( .A(n226), .B(n48), .Z(n49) );
  OR2 C75 ( .A(n437), .B(n69), .Z(n52) );
  OR2 C80 ( .A(n446), .B(n32), .Z(n55) );
  OR2 C83 ( .A(n223), .B(n455), .Z(n58) );
  OR2 C84 ( .A(n224), .B(n58), .Z(n59) );
  OR2 C85 ( .A(n225), .B(n59), .Z(n60) );
  OR2 C88 ( .A(n454), .B(n222), .Z(n63) );
  OR2 C89 ( .A(n224), .B(n63), .Z(n64) );
  OR2 C90 ( .A(n225), .B(n64), .Z(n65) );
  OR2 C941 ( .A(n453), .B(n31), .Z(n68) );
  OR2 C951 ( .A(n225), .B(n68), .Z(n69) );
  OR2 C100 ( .A(n454), .B(n455), .Z(n71) );
  OR2 C101 ( .A(n453), .B(n71), .Z(n72) );
  OR2 C1021 ( .A(n225), .B(n72), .Z(n73) );
  OR2 C1031 ( .A(n226), .B(n73), .Z(n74) );
  OR2 C1081 ( .A(n226), .B(n33), .Z(n76) );
  OR2 C1141 ( .A(n226), .B(n60), .Z(n78) );
  OR2 C120 ( .A(n226), .B(n65), .Z(n80) );
  OR2 C126 ( .A(n226), .B(n69), .Z(n82) );
  OR2 C1321 ( .A(n226), .B(n55), .Z(n84) );
  OR2 C140 ( .A(n446), .B(n72), .Z(n86) );
  OR2 C141 ( .A(n226), .B(n86), .Z(n87) );
  OR2 C148 ( .A(n437), .B(n55), .Z(n89) );
  OR2 C154 ( .A(n437), .B(n33), .Z(n91) );
  AN2 C159 ( .A(n226), .B(n30), .Z(n93) );
  OR2 C167 ( .A(n437), .B(n73), .Z(n94) );
  OR2 C174 ( .A(n224), .B(n71), .Z(n96) );
  OR2 C175 ( .A(n446), .B(n96), .Z(n97) );
  OR2 C176 ( .A(n437), .B(n97), .Z(n98) );
  OR2 C183 ( .A(n453), .B(n58), .Z(n100) );
  OR2 C184 ( .A(n446), .B(n100), .Z(n101) );
  OR2 C185 ( .A(n437), .B(n101), .Z(n102) );
  OR2 C192 ( .A(n453), .B(n63), .Z(n104) );
  OR2 C193 ( .A(n446), .B(n104), .Z(n105) );
  OR2 C194 ( .A(n437), .B(n105), .Z(n106) );
  OR2 C202 ( .A(n437), .B(n48), .Z(n108) );
  OR2 C206 ( .A(n111), .B(n451), .Z(n[5]) );
  AN2 C207 ( .A(n223), .B(n452), .Z(n111) );
  OR2 C209 ( .A(n112), .B(n435), .Z(n[6]) );
  OR2 C210 ( .A(n224), .B(n451), .Z(n112) );
  AN2 C211 ( .A(n225), .B(n452), .Z(n[7]) );
  OR2 C213 ( .A(n113), .B(n115), .Z(n[8]) );
  OR2 C215 ( .A(n114), .B(n447), .Z(n115) );
  OR2 C216 ( .A(n449), .B(n448), .Z(n114) );
  OR2 C217 ( .A(n125), .B(n126), .Z(n[9]) );
  OR2 C218 ( .A(n124), .B(n93), .Z(n125) );
  OR2 C219 ( .A(n123), .B(n436), .Z(n124) );
  OR2 C220 ( .A(n122), .B(n445), .Z(n123) );
  OR2 C221 ( .A(n117), .B(n121), .Z(n122) );
  AN2 C222 ( .A(n450), .B(n116), .Z(n117) );
  AN2 C224 ( .A(n120), .B(n437), .Z(n121) );
  AN2 C225 ( .A(n118), .B(n119), .Z(n120) );
  AN2 C229 ( .A(n429), .B(n221), .Z(n126) );
  OR2 C230 ( .A(n131), .B(n435), .Z(n10) );
  OR2 C231 ( .A(n130), .B(n438), .Z(n131) );
  OR2 C232 ( .A(n129), .B(n439), .Z(n130) );
  OR2 C233 ( .A(n128), .B(n440), .Z(n129) );
  OR2 C234 ( .A(n127), .B(n441), .Z(n128) );
  OR2 C235 ( .A(n443), .B(n442), .Z(n127) );
  OR2 C236 ( .A(n136), .B(n137), .Z(n11) );
  OR2 C237 ( .A(n135), .B(n93), .Z(n136) );
  OR2 C238 ( .A(n134), .B(n430), .Z(n135) );
  OR2 C239 ( .A(n133), .B(n431), .Z(n134) );
  OR2 C240 ( .A(n132), .B(n432), .Z(n133) );
  OR2 C241 ( .A(n434), .B(n433), .Z(n132) );
  AN2 C242 ( .A(n429), .B(n221), .Z(n137) );
  AN2 C243 ( .A(n142), .B(n36), .Z(n13) );
  OR2 C244 ( .A(n141), .B(n221), .Z(n142) );
  OR2 C245 ( .A(n138), .B(n140), .Z(n141) );
  AN2 C246 ( .A(n419), .B(n418), .Z(n138) );
  AN2 C247 ( .A(n460), .B(n39), .Z(n140) );
  AN2 C249 ( .A(n227), .B(n417), .Z(n14) );
  OR2 C251 ( .A(n228), .B(n424), .Z(n15) );
  OR2 C252 ( .A(n145), .B(n13), .Z(n16) );
  AN2 C253 ( .A(n147), .B(n423), .Z(n145) );
  OR2 C256 ( .A(n424), .B(n422), .Z(n17) );
  AN2 C257 ( .A(n146), .B(n147), .Z(n18) );
  AN2 C258 ( .A(n429), .B(n221), .Z(n146) );
  OR2 C260 ( .A(n150), .B(n429), .Z(n19) );
  OR2 C261 ( .A(n149), .B(n430), .Z(n150) );
  OR2 C262 ( .A(n148), .B(n431), .Z(n149) );
  OR2 C263 ( .A(n433), .B(n432), .Z(n148) );
  OR2 C265 ( .A(n10), .B(n11), .Z(n151) );
  AN2 C266 ( .A(n219), .B(n154), .Z(n4) );
  OR2 C269 ( .A(n17), .B(n36), .Z(n153) );
  AN2 C270 ( .A(n421), .B(n3), .Z(n20) );
  OR2 C272 ( .A(n160), .B(n162), .Z(n21) );
  OR2 C273 ( .A(n157), .B(n159), .Z(n160) );
  AN2 C274 ( .A(n420), .B(n10), .Z(n157) );
  AN2 C276 ( .A(n20), .B(n158), .Z(n159) );
  OR2 C277 ( .A(n444), .B(n11), .Z(n158) );
  AN2 C278 ( .A(n428), .B(n221), .Z(n162) );
  OR2 C280 ( .A(n164), .B(n166), .Z(n22) );
  AN2 C281 ( .A(n460), .B(n163), .Z(n164) );
  OR2 C283 ( .A(n17), .B(n18), .Z(n163) );
  AN2 C284 ( .A(n419), .B(n165), .Z(n166) );
  OR2 C285 ( .A(n425), .B(n36), .Z(n165) );
  AN2 C136 ( .A(TXDATAK), .B(n175), .Z(n171) );
  AN2 C135 ( .A(n193), .B(n185), .Z(n172) );
  OR2 C134 ( .A(n172), .B(n171), .Z(n170) );
  AN2 C133 ( .A(n170), .B(CNTL_RESETN_P0), .Z(n169) );
  AN2 C132 ( .A(n169), .B(n206), .Z(n168) );
  AN2 C131 ( .A(n168), .B(n173), .Z(n167) );
  AN2 C130 ( .A(n167), .B(CNTL_TXEnable_P0), .Z(assertion_shengyushen) );
  IV I_11 ( .A(CNTL_Loopback_P0), .Z(n206) );
  AN2 C119 ( .A(CNTL_TXEnable_P0), .B(n173), .Z(U6_DATA2_0) );
  IV I_9 ( .A(TXELECIDLE), .Z(n173) );
  AN2 C117 ( .A(RST_BeaconEnable_R0), .B(n173), .Z(HSS_TXBEACONCMD) );
  IV I_8 ( .A(CNTL_RESETN_P0), .Z(n174) );
  IV I_7 ( .A(n176), .Z(n175) );
  OR2 C108 ( .A(TXDATA[0]), .B(n177), .Z(n176) );
  OR2 C107 ( .A(TXDATA[1]), .B(n178), .Z(n177) );
  OR2 C106 ( .A(n183), .B(n179), .Z(n178) );
  OR2 C105 ( .A(n190), .B(n180), .Z(n179) );
  OR2 C104 ( .A(n184), .B(n181), .Z(n180) );
  OR2 C103 ( .A(n191), .B(n182), .Z(n181) );
  OR2 C102 ( .A(TXDATA[6]), .B(TXDATA[7]), .Z(n182) );
  IV I_6 ( .A(TXDATA[2]), .Z(n183) );
  IV I_5 ( .A(TXDATA[4]), .Z(n184) );
  IV I_4 ( .A(n186), .Z(n185) );
  OR2 C96 ( .A(n190), .B(n187), .Z(n186) );
  OR2 C95 ( .A(TXDATA[4]), .B(n188), .Z(n187) );
  OR2 C94 ( .A(n191), .B(n189), .Z(n188) );
  OR2 C93 ( .A(n192), .B(TXDATA[7]), .Z(n189) );
  IV I_3 ( .A(TXDATA[3]), .Z(n190) );
  IV I_2 ( .A(TXDATA[5]), .Z(n191) );
  IV I_1 ( .A(TXDATA[6]), .Z(n192) );
  IV I_0 ( .A(TXDATAK), .Z(n193) );
  FD1 InputDataK_P0_reg ( .D(n416), .CP(PCLK250), .Q(n221) );
  FD1 InputCompliance_P0_reg ( .D(n415), .CP(PCLK250), .Q(n220) );
  FD1 InputData_P0_reg_7_ ( .D(n414), .CP(PCLK250), .Q(n229) );
  FD1 InputData_P0_reg_6_ ( .D(n413), .CP(PCLK250), .Q(n228) );
  FD1 InputData_P0_reg_5_ ( .D(n412), .CP(PCLK250), .Q(n227) );
  FD1 InputData_P0_reg_4_ ( .D(n411), .CP(PCLK250), .Q(n226) );
  FD1 InputData_P0_reg_3_ ( .D(n410), .CP(PCLK250), .Q(n225) );
  FD1 InputData_P0_reg_2_ ( .D(n409), .CP(PCLK250), .Q(n224) );
  FD1 InputData_P0_reg_1_ ( .D(n408), .CP(PCLK250), .Q(n223) );
  FD1 InputData_P0_reg_0_ ( .D(n407), .CP(PCLK250), .Q(n222) );
  FD1 InputDataEnable_P0_reg ( .D(U6_Z_0), .CP(PCLK250), .Q(n219) );
  FD1 OutputElecIdle_P0_reg ( .D(U4_Z_0), .CP(PCLK250), .Q(HSS_TXELECIDLE) );
  FD1 DISPARITY_P0_reg ( .D(n4), .CP(PCLK250), .Q(n3) );
  FD1 OutputData_P0_reg_7_ ( .D(n406), .CP(PCLK250), .Q(HSS_TXD[7]) );
  FD1 OutputData_P0_reg_8_ ( .D(n405), .CP(PCLK250), .Q(HSS_TXD[8]) );
  FD1 OutputData_P0_reg_4_ ( .D(n404), .CP(PCLK250), .Q(HSS_TXD[4]) );
  FD1 OutputData_P0_reg_9_ ( .D(n403), .CP(PCLK250), .Q(HSS_TXD[9]) );
  FD1 OutputData_P0_reg_6_ ( .D(n402), .CP(PCLK250), .Q(HSS_TXD[6]) );
  FD1 OutputData_P0_reg_5_ ( .D(n401), .CP(PCLK250), .Q(HSS_TXD[5]) );
  FD1 OutputData_P0_reg_0_ ( .D(n400), .CP(PCLK250), .Q(HSS_TXD[0]) );
  FD1 OutputData_P0_reg_1_ ( .D(n399), .CP(PCLK250), .Q(HSS_TXD[1]) );
  FD1 OutputData_P0_reg_2_ ( .D(n398), .CP(PCLK250), .Q(HSS_TXD[2]) );
  FD1 OutputData_P0_reg_3_ ( .D(n397), .CP(PCLK250), .Q(HSS_TXD[3]) );
  AN2 U88 ( .A(U6_DATA2_0), .B(TXDATA[0]), .Z(n351) );
  AN2 U91 ( .A(TXDATA[1]), .B(U6_DATA2_0), .Z(n354) );
  AN2 U94 ( .A(TXDATA[2]), .B(U6_DATA2_0), .Z(n356) );
  AN2 U97 ( .A(TXDATA[3]), .B(U6_DATA2_0), .Z(n358) );
  AN2 U100 ( .A(TXDATA[4]), .B(U6_DATA2_0), .Z(n360) );
  AN2 U103 ( .A(TXDATA[5]), .B(U6_DATA2_0), .Z(n362) );
  AN2 U106 ( .A(TXDATA[6]), .B(U6_DATA2_0), .Z(n364) );
  AN2 U109 ( .A(TXDATA[7]), .B(U6_DATA2_0), .Z(n366) );
  AN2 U112 ( .A(TXCOMPLIANCE), .B(U6_DATA2_0), .Z(n368) );
  IV U115 ( .A(U6_DATA2_0), .Z(n353) );
  AN2 U116 ( .A(TXDATAK), .B(U6_DATA2_0), .Z(n370) );
  AN2 U181 ( .A(CNTL_RESETN_P0), .B(U6_DATA2_0), .Z(U6_Z_0) );
  IV U194 ( .A(n30), .Z(n452) );
  IV U195 ( .A(n33), .Z(n451) );
  IV U196 ( .A(n46), .Z(n450) );
  IV U197 ( .A(n60), .Z(n449) );
  IV U198 ( .A(n65), .Z(n448) );
  IV U199 ( .A(n69), .Z(n447) );
  IV U200 ( .A(n49), .Z(n445) );
  IV U201 ( .A(n74), .Z(n444) );
  IV U202 ( .A(n76), .Z(n443) );
  IV U203 ( .A(n78), .Z(n442) );
  IV U204 ( .A(n80), .Z(n441) );
  IV U205 ( .A(n82), .Z(n440) );
  IV U206 ( .A(n84), .Z(n439) );
  IV U207 ( .A(n87), .Z(n438) );
  IV U208 ( .A(n52), .Z(n436) );
  IV U209 ( .A(n89), .Z(n435) );
  IV U210 ( .A(n91), .Z(n434) );
  IV U211 ( .A(n94), .Z(n433) );
  IV U212 ( .A(n98), .Z(n432) );
  IV U213 ( .A(n102), .Z(n431) );
  IV U214 ( .A(n106), .Z(n430) );
  IV U215 ( .A(n108), .Z(n429) );
  IV U216 ( .A(n19), .Z(n428) );
  IV U217 ( .A(n26), .Z(n425) );
  IV U218 ( .A(n41), .Z(n424) );
  IV U219 ( .A(n44), .Z(n422) );
  IV U220 ( .A(n220), .Z(n421) );
  IV U221 ( .A(n37), .Z(n418) );
  IV U222 ( .A(n13), .Z(n417) );
  OR2 U223 ( .A(n461), .B(n370), .Z(n416) );
  AN2 U224 ( .A(n353), .B(n221), .Z(n461) );
  OR2 U225 ( .A(n462), .B(n368), .Z(n415) );
  AN2 U226 ( .A(n353), .B(n220), .Z(n462) );
  OR2 U227 ( .A(n463), .B(n366), .Z(n414) );
  AN2 U228 ( .A(n353), .B(n229), .Z(n463) );
  OR2 U229 ( .A(n464), .B(n364), .Z(n413) );
  AN2 U230 ( .A(n353), .B(n228), .Z(n464) );
  OR2 U231 ( .A(n465), .B(n362), .Z(n412) );
  AN2 U232 ( .A(n353), .B(n227), .Z(n465) );
  OR2 U233 ( .A(n466), .B(n360), .Z(n411) );
  AN2 U234 ( .A(n353), .B(n226), .Z(n466) );
  OR2 U235 ( .A(n467), .B(n358), .Z(n410) );
  AN2 U236 ( .A(n353), .B(n225), .Z(n467) );
  OR2 U237 ( .A(n468), .B(n356), .Z(n409) );
  AN2 U238 ( .A(n353), .B(n224), .Z(n468) );
  OR2 U239 ( .A(n469), .B(n354), .Z(n408) );
  AN2 U240 ( .A(n353), .B(n223), .Z(n469) );
  OR2 U241 ( .A(n470), .B(n351), .Z(n407) );
  AN2 U242 ( .A(n353), .B(n222), .Z(n470) );
  OR2 U243 ( .A(n471), .B(n472), .Z(n406) );
  OR2 U244 ( .A(n473), .B(n474), .Z(n472) );
  AN2 U245 ( .A(HSS_TXD[7]), .B(n475), .Z(n474) );
  AN2 U246 ( .A(RX_LoopbackData_P2[7]), .B(n476), .Z(n473) );
  OR2 U247 ( .A(n477), .B(n478), .Z(n471) );
  AN2 U248 ( .A(n479), .B(n15), .Z(n478) );
  AN2 U249 ( .A(n480), .B(n481), .Z(n477) );
  IV U250 ( .A(n15), .Z(n481) );
  OR2 U251 ( .A(n482), .B(n483), .Z(n405) );
  OR2 U252 ( .A(n484), .B(n485), .Z(n483) );
  AN2 U253 ( .A(HSS_TXD[8]), .B(n475), .Z(n485) );
  AN2 U254 ( .A(RX_LoopbackData_P2[8]), .B(n476), .Z(n484) );
  OR2 U255 ( .A(n486), .B(n487), .Z(n482) );
  AN2 U256 ( .A(n479), .B(n229), .Z(n487) );
  AN2 U257 ( .A(n480), .B(n423), .Z(n486) );
  IV U258 ( .A(n229), .Z(n423) );
  OR2 U259 ( .A(n488), .B(n489), .Z(n404) );
  OR2 U260 ( .A(n490), .B(n491), .Z(n489) );
  AN2 U261 ( .A(RX_LoopbackData_P2[4]), .B(n476), .Z(n491) );
  AN2 U262 ( .A(n492), .B(U5_DATA2_4), .Z(n490) );
  AN2 U263 ( .A(HSS_TXD[4]), .B(n475), .Z(n488) );
  OR2 U264 ( .A(n493), .B(n494), .Z(n403) );
  OR2 U265 ( .A(n495), .B(n496), .Z(n494) );
  AN2 U266 ( .A(HSS_TXD[9]), .B(n475), .Z(n496) );
  AN2 U267 ( .A(RX_LoopbackData_P2[9]), .B(n476), .Z(n495) );
  OR2 U268 ( .A(n497), .B(n498), .Z(n493) );
  AN2 U269 ( .A(n16), .B(n479), .Z(n498) );
  AN2 U270 ( .A(n480), .B(n499), .Z(n497) );
  IV U271 ( .A(n16), .Z(n499) );
  OR2 U272 ( .A(n500), .B(n501), .Z(n402) );
  OR2 U273 ( .A(n502), .B(n503), .Z(n501) );
  AN2 U274 ( .A(HSS_TXD[6]), .B(n475), .Z(n503) );
  AN2 U275 ( .A(RX_LoopbackData_P2[6]), .B(n476), .Z(n502) );
  OR2 U276 ( .A(n504), .B(n505), .Z(n500) );
  AN2 U277 ( .A(n14), .B(n479), .Z(n505) );
  AN2 U278 ( .A(n506), .B(n492), .Z(n479) );
  IV U279 ( .A(n22), .Z(n506) );
  AN2 U280 ( .A(n480), .B(n507), .Z(n504) );
  IV U281 ( .A(n14), .Z(n507) );
  AN2 U282 ( .A(n492), .B(n22), .Z(n480) );
  OR2 U283 ( .A(n508), .B(n509), .Z(n401) );
  OR2 U284 ( .A(n510), .B(n511), .Z(n509) );
  AN2 U285 ( .A(RX_LoopbackData_P2[5]), .B(n476), .Z(n511) );
  AN2 U286 ( .A(n492), .B(U5_DATA2_5), .Z(n510) );
  AN2 U287 ( .A(HSS_TXD[5]), .B(n475), .Z(n508) );
  OR2 U288 ( .A(n512), .B(n513), .Z(n400) );
  OR2 U289 ( .A(n514), .B(n515), .Z(n513) );
  AN2 U290 ( .A(HSS_TXD[0]), .B(n475), .Z(n515) );
  AN2 U291 ( .A(RX_LoopbackData_P2[0]), .B(n476), .Z(n514) );
  OR2 U292 ( .A(n516), .B(n517), .Z(n512) );
  AN2 U293 ( .A(n518), .B(n222), .Z(n517) );
  AN2 U294 ( .A(n519), .B(n455), .Z(n516) );
  OR2 U295 ( .A(n520), .B(n521), .Z(n399) );
  OR2 U296 ( .A(n522), .B(n523), .Z(n521) );
  AN2 U297 ( .A(HSS_TXD[1]), .B(n475), .Z(n523) );
  AN2 U298 ( .A(RX_LoopbackData_P2[1]), .B(n476), .Z(n522) );
  OR2 U299 ( .A(n524), .B(n525), .Z(n520) );
  AN2 U300 ( .A(n[5]), .B(n518), .Z(n525) );
  AN2 U301 ( .A(n519), .B(n526), .Z(n524) );
  IV U302 ( .A(n[5]), .Z(n526) );
  OR2 U303 ( .A(n527), .B(n528), .Z(n398) );
  OR2 U304 ( .A(n529), .B(n530), .Z(n528) );
  AN2 U305 ( .A(HSS_TXD[2]), .B(n475), .Z(n530) );
  AN2 U306 ( .A(RX_LoopbackData_P2[2]), .B(n476), .Z(n529) );
  OR2 U307 ( .A(n531), .B(n532), .Z(n527) );
  AN2 U308 ( .A(n[6]), .B(n518), .Z(n532) );
  AN2 U309 ( .A(n519), .B(n533), .Z(n531) );
  IV U310 ( .A(n[6]), .Z(n533) );
  OR2 U311 ( .A(n534), .B(n535), .Z(n397) );
  OR2 U312 ( .A(n536), .B(n537), .Z(n535) );
  AN2 U313 ( .A(HSS_TXD[3]), .B(n475), .Z(n537) );
  AN2 U314 ( .A(RX_LoopbackData_P2[3]), .B(n476), .Z(n536) );
  AN2 U315 ( .A(n219), .B(CNTL_Loopback_P0), .Z(n476) );
  OR2 U316 ( .A(n538), .B(n539), .Z(n534) );
  AN2 U317 ( .A(n[7]), .B(n518), .Z(n539) );
  AN2 U318 ( .A(n540), .B(n492), .Z(n518) );
  AN2 U319 ( .A(n519), .B(n541), .Z(n538) );
  IV U320 ( .A(n[7]), .Z(n541) );
  AN2 U321 ( .A(n492), .B(n21), .Z(n519) );
  AN2 U322 ( .A(n206), .B(n219), .Z(n492) );
  OR2 U323 ( .A(n542), .B(n543), .Z(n154) );
  IV U324 ( .A(n544), .Z(n543) );
  OR2 U325 ( .A(n460), .B(n153), .Z(n544) );
  AN2 U326 ( .A(n153), .B(n460), .Z(n542) );
  IV U327 ( .A(n419), .Z(n460) );
  OR2 U328 ( .A(n545), .B(n546), .Z(n419) );
  AN2 U329 ( .A(n151), .B(n420), .Z(n546) );
  IV U330 ( .A(n547), .Z(n545) );
  OR2 U331 ( .A(n420), .B(n151), .Z(n547) );
  IV U332 ( .A(n20), .Z(n420) );
  OR2 U333 ( .A(n548), .B(n549), .Z(n147) );
  AN2 U334 ( .A(n227), .B(n426), .Z(n549) );
  IV U335 ( .A(n228), .Z(n426) );
  AN2 U336 ( .A(n228), .B(n427), .Z(n548) );
  IV U337 ( .A(n227), .Z(n427) );
  OR2 U338 ( .A(n550), .B(n551), .Z(n119) );
  AN2 U339 ( .A(n224), .B(n446), .Z(n551) );
  IV U340 ( .A(n225), .Z(n446) );
  AN2 U341 ( .A(n225), .B(n453), .Z(n550) );
  IV U342 ( .A(n224), .Z(n453) );
  OR2 U343 ( .A(n552), .B(n553), .Z(n118) );
  AN2 U344 ( .A(n222), .B(n454), .Z(n553) );
  IV U345 ( .A(n223), .Z(n454) );
  AN2 U346 ( .A(n223), .B(n455), .Z(n552) );
  IV U347 ( .A(n222), .Z(n455) );
  OR2 U348 ( .A(n554), .B(n555), .Z(n116) );
  IV U349 ( .A(n556), .Z(n555) );
  OR2 U350 ( .A(n437), .B(n28), .Z(n556) );
  AN2 U351 ( .A(n28), .B(n437), .Z(n554) );
  AN2 U352 ( .A(n557), .B(n558), .Z(n113) );
  IV U353 ( .A(n559), .Z(n558) );
  AN2 U354 ( .A(n437), .B(n55), .Z(n559) );
  OR2 U355 ( .A(n55), .B(n437), .Z(n557) );
  IV U356 ( .A(n226), .Z(n437) );
  OR2 U357 ( .A(n560), .B(n561), .Z(U5_DATA2_5) );
  IV U358 ( .A(n562), .Z(n561) );
  OR2 U359 ( .A(n540), .B(n[9]), .Z(n562) );
  AN2 U360 ( .A(n[9]), .B(n540), .Z(n560) );
  OR2 U361 ( .A(n563), .B(n564), .Z(U5_DATA2_4) );
  IV U362 ( .A(n565), .Z(n564) );
  OR2 U363 ( .A(n540), .B(n[8]), .Z(n565) );
  AN2 U364 ( .A(n[8]), .B(n540), .Z(n563) );
  IV U365 ( .A(n21), .Z(n540) );
  OR2 U366 ( .A(n566), .B(n174), .Z(U4_Z_0) );
  AN2 U367 ( .A(CNTL_RESETN_P0), .B(n475), .Z(n566) );
  IV U368 ( .A(n219), .Z(n475) );
endmodule

