
module PCIEXP_TX ( PCLK250, RST_BeaconEnable_R0, CNTL_RESETN_P0, 
        CNTL_Loopback_P0, CNTL_TXEnable_P0, RX_LoopbackData_P2, TXCOMPLIANCE, 
        TXDATA, TXDATAK, TXELECIDLE, HSS_TXBEACONCMD, HSS_TXD, HSS_TXELECIDLE, 
        assertion_shengyushen );
  input [9:0] RX_LoopbackData_P2;
  input [7:0] TXDATA;
  output [9:0] HSS_TXD;
  input PCLK250, RST_BeaconEnable_R0, CNTL_RESETN_P0, CNTL_Loopback_P0,
         CNTL_TXEnable_P0, TXCOMPLIANCE, TXDATAK, TXELECIDLE;
  output HSS_TXBEACONCMD, HSS_TXELECIDLE, assertion_shengyushen;
  wire   n4, n5, n11, n12, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n38, n39, n41, n42, n43, n44, n45, n46, n47, n48, n50, n52,
         n53, n54, n57, n60, n61, n62, n63, n64, n65, n66, n69, n70, n72, n74,
         n75, n78, n81, n83, n84, n85, n87, n88, n89, n92, n93, n95, n96, n97,
         n98, n100, n102, n104, n106, n108, n110, n111, n113, n115, n117, n118,
         n120, n121, n122, n124, n125, n126, n128, n129, n130, n132, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n164, n165, n166, n169, n170, n171,
         n172, n173, n174, n175, n177, n178, n181, n182, n183, n184, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         U7_Z_0, U7_DATA2_0, U5_Z_0, U4_DATA2_4, U4_DATA2_5, n399, n446, n448,
         n449, n451, n453, n455, n457, n459, n461, n463, n465, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666;
  wire   [6:10] n;

  OR2 C52 ( .A(n523), .B(n524), .Z(n38) );
  OR2 C53 ( .A(n320), .B(n38), .Z(n39) );
  AN2 C55 ( .A(n319), .B(n318), .Z(n41) );
  AN2 C56 ( .A(n320), .B(n41), .Z(n42) );
  AN2 C57 ( .A(n314), .B(n313), .Z(n43) );
  AN2 C58 ( .A(n315), .B(n43), .Z(n44) );
  AN2 C59 ( .A(n316), .B(n44), .Z(n45) );
  OR2 C60 ( .A(n314), .B(n313), .Z(n46) );
  OR2 C61 ( .A(n315), .B(n46), .Z(n47) );
  OR2 C62 ( .A(n316), .B(n47), .Z(n48) );
  OR2 C64 ( .A(U4_DATA2_5), .B(U4_DATA2_4), .Z(n50) );
  AN2 C66 ( .A(U4_DATA2_5), .B(U4_DATA2_4), .Z(n52) );
  OR2 C69 ( .A(n319), .B(n318), .Z(n53) );
  OR2 C70 ( .A(n320), .B(n53), .Z(n54) );
  OR2 C74 ( .A(n518), .B(n53), .Z(n57) );
  OR2 C77 ( .A(n319), .B(n320), .Z(n60) );
  OR2 C78 ( .A(n318), .B(n60), .Z(n61) );
  OR2 C79 ( .A(n317), .B(n61), .Z(n62) );
  OR2 C80 ( .A(n316), .B(n62), .Z(n63) );
  OR2 C81 ( .A(n315), .B(n63), .Z(n64) );
  OR2 C82 ( .A(n314), .B(n64), .Z(n65) );
  OR2 C83 ( .A(n552), .B(n65), .Z(n66) );
  OR2 C91 ( .A(n551), .B(n64), .Z(n69) );
  OR2 C92 ( .A(n313), .B(n69), .Z(n70) );
  OR2 C94 ( .A(n316), .B(n315), .Z(n72) );
  OR2 C1011 ( .A(n543), .B(n92), .Z(n74) );
  OR2 C1021 ( .A(n317), .B(n74), .Z(n75) );
  OR2 C109 ( .A(n534), .B(n93), .Z(n78) );
  OR2 C1141 ( .A(n543), .B(n47), .Z(n81) );
  OR2 C117 ( .A(n314), .B(n552), .Z(n83) );
  OR2 C118 ( .A(n315), .B(n83), .Z(n84) );
  OR2 C119 ( .A(n316), .B(n84), .Z(n85) );
  OR2 C1221 ( .A(n551), .B(n313), .Z(n87) );
  OR2 C1231 ( .A(n315), .B(n87), .Z(n88) );
  OR2 C1241 ( .A(n316), .B(n88), .Z(n89) );
  OR2 C1281 ( .A(n550), .B(n46), .Z(n92) );
  OR2 C129 ( .A(n316), .B(n92), .Z(n93) );
  OR2 C1341 ( .A(n551), .B(n552), .Z(n95) );
  OR2 C1351 ( .A(n550), .B(n95), .Z(n96) );
  OR2 C1361 ( .A(n316), .B(n96), .Z(n97) );
  OR2 C1371 ( .A(n317), .B(n97), .Z(n98) );
  OR2 C142 ( .A(n317), .B(n48), .Z(n100) );
  OR2 C1481 ( .A(n317), .B(n85), .Z(n102) );
  OR2 C154 ( .A(n317), .B(n89), .Z(n104) );
  OR2 C1601 ( .A(n317), .B(n93), .Z(n106) );
  OR2 C1661 ( .A(n317), .B(n81), .Z(n108) );
  OR2 C174 ( .A(n543), .B(n96), .Z(n110) );
  OR2 C1751 ( .A(n317), .B(n110), .Z(n111) );
  OR2 C182 ( .A(n534), .B(n81), .Z(n113) );
  OR2 C188 ( .A(n534), .B(n48), .Z(n115) );
  AN2 C1931 ( .A(n317), .B(n45), .Z(n117) );
  OR2 C201 ( .A(n534), .B(n97), .Z(n118) );
  OR2 C2081 ( .A(n315), .B(n95), .Z(n120) );
  OR2 C2091 ( .A(n543), .B(n120), .Z(n121) );
  OR2 C2101 ( .A(n534), .B(n121), .Z(n122) );
  OR2 C217 ( .A(n550), .B(n83), .Z(n124) );
  OR2 C218 ( .A(n543), .B(n124), .Z(n125) );
  OR2 C219 ( .A(n534), .B(n125), .Z(n126) );
  OR2 C226 ( .A(n550), .B(n87), .Z(n128) );
  OR2 C227 ( .A(n543), .B(n128), .Z(n129) );
  OR2 C228 ( .A(n534), .B(n129), .Z(n130) );
  OR2 C236 ( .A(n534), .B(n74), .Z(n132) );
  OR2 C241 ( .A(n135), .B(n548), .Z(n[6]) );
  AN2 C242 ( .A(n314), .B(n549), .Z(n135) );
  OR2 C244 ( .A(n136), .B(n532), .Z(n[7]) );
  OR2 C245 ( .A(n315), .B(n548), .Z(n136) );
  AN2 C2461 ( .A(n316), .B(n549), .Z(n[8]) );
  OR2 C2481 ( .A(n137), .B(n139), .Z(n[9]) );
  OR2 C250 ( .A(n138), .B(n544), .Z(n139) );
  OR2 C2511 ( .A(n546), .B(n545), .Z(n138) );
  OR2 C252 ( .A(n149), .B(n150), .Z(n[10]) );
  OR2 C2531 ( .A(n148), .B(n117), .Z(n149) );
  OR2 C254 ( .A(n147), .B(n533), .Z(n148) );
  OR2 C255 ( .A(n146), .B(n542), .Z(n147) );
  OR2 C256 ( .A(n141), .B(n145), .Z(n146) );
  AN2 C257 ( .A(n547), .B(n140), .Z(n141) );
  AN2 C259 ( .A(n144), .B(n534), .Z(n145) );
  AN2 C260 ( .A(n142), .B(n143), .Z(n144) );
  AN2 C2641 ( .A(n526), .B(n312), .Z(n150) );
  OR2 C2651 ( .A(n155), .B(n532), .Z(n11) );
  OR2 C2661 ( .A(n154), .B(n535), .Z(n155) );
  OR2 C2671 ( .A(n153), .B(n536), .Z(n154) );
  OR2 C2681 ( .A(n152), .B(n537), .Z(n153) );
  OR2 C2691 ( .A(n151), .B(n538), .Z(n152) );
  OR2 C2701 ( .A(n540), .B(n539), .Z(n151) );
  OR2 C2711 ( .A(n160), .B(n161), .Z(n12) );
  OR2 C2721 ( .A(n159), .B(n117), .Z(n160) );
  OR2 C2731 ( .A(n158), .B(n527), .Z(n159) );
  OR2 C2741 ( .A(n157), .B(n528), .Z(n158) );
  OR2 C2751 ( .A(n156), .B(n529), .Z(n157) );
  OR2 C2761 ( .A(n531), .B(n530), .Z(n156) );
  AN2 C2771 ( .A(n526), .B(n312), .Z(n161) );
  AN2 C2781 ( .A(n166), .B(n42), .Z(n24) );
  OR2 C2791 ( .A(n165), .B(n312), .Z(n166) );
  OR2 C2801 ( .A(n162), .B(n164), .Z(n165) );
  AN2 C281 ( .A(n23), .B(n513), .Z(n162) );
  AN2 C282 ( .A(n514), .B(n52), .Z(n164) );
  AN2 C284 ( .A(n318), .B(n512), .Z(n25) );
  OR2 C286 ( .A(n319), .B(n521), .Z(n26) );
  OR2 C287 ( .A(n169), .B(n24), .Z(n27) );
  AN2 C288 ( .A(n171), .B(n518), .Z(n169) );
  OR2 C291 ( .A(n521), .B(n517), .Z(n28) );
  AN2 C292 ( .A(n170), .B(n171), .Z(n29) );
  AN2 C293 ( .A(n526), .B(n312), .Z(n170) );
  OR2 C295 ( .A(n174), .B(n526), .Z(n30) );
  OR2 C296 ( .A(n173), .B(n527), .Z(n174) );
  OR2 C297 ( .A(n172), .B(n528), .Z(n173) );
  OR2 C298 ( .A(n530), .B(n529), .Z(n172) );
  OR2 C300 ( .A(n11), .B(n12), .Z(n175) );
  AN2 C301 ( .A(n310), .B(n178), .Z(n5) );
  OR2 C304 ( .A(n28), .B(n42), .Z(n177) );
  AN2 C305 ( .A(n516), .B(n4), .Z(n31) );
  OR2 C307 ( .A(n184), .B(n186), .Z(n32) );
  OR2 C308 ( .A(n181), .B(n183), .Z(n184) );
  AN2 C309 ( .A(n515), .B(n11), .Z(n181) );
  AN2 C311 ( .A(n31), .B(n182), .Z(n183) );
  OR2 C312 ( .A(n541), .B(n12), .Z(n182) );
  AN2 C313 ( .A(n525), .B(n312), .Z(n186) );
  OR2 C315 ( .A(n188), .B(n190), .Z(n33) );
  AN2 C316 ( .A(n514), .B(n187), .Z(n188) );
  OR2 C318 ( .A(n28), .B(n29), .Z(n187) );
  AN2 C319 ( .A(n23), .B(n189), .Z(n190) );
  OR2 C320 ( .A(n522), .B(n42), .Z(n189) );
  OR2 C331 ( .A(n520), .B(n519), .Z(n34) );
  OR2 C280 ( .A(n274), .B(n266), .Z(n206) );
  OR2 C279 ( .A(n206), .B(n257), .Z(n205) );
  OR2 C278 ( .A(n205), .B(n248), .Z(n204) );
  OR2 C277 ( .A(n204), .B(n241), .Z(n203) );
  OR2 C276 ( .A(n203), .B(n233), .Z(n202) );
  OR2 C275 ( .A(n202), .B(n226), .Z(n201) );
  OR2 C274 ( .A(n201), .B(n219), .Z(n200) );
  OR2 C273 ( .A(n200), .B(n215), .Z(n199) );
  OR2 C272 ( .A(n199), .B(n213), .Z(n198) );
  OR2 C271 ( .A(n198), .B(n210), .Z(n197) );
  AN2 C270 ( .A(TXDATAK), .B(n197), .Z(n196) );
  OR2 C269 ( .A(n285), .B(n196), .Z(n195) );
  AN2 C268 ( .A(n195), .B(CNTL_RESETN_P0), .Z(n194) );
  AN2 C267 ( .A(n194), .B(CNTL_TXEnable_P0), .Z(n193) );
  AN2 C266 ( .A(n193), .B(n209), .Z(n192) );
  AN2 C265 ( .A(n192), .B(n208), .Z(n191) );
  AN2 C264 ( .A(n191), .B(TXCOMPLIANCE), .Z(assertion_shengyushen) );
  AN2 C253 ( .A(CNTL_TXEnable_P0), .B(n209), .Z(U7_DATA2_0) );
  AN2 C251 ( .A(RST_BeaconEnable_R0), .B(n209), .Z(HSS_TXBEACONCMD) );
  IV I_22 ( .A(CNTL_RESETN_P0), .Z(n207) );
  IV I_21 ( .A(CNTL_Loopback_P0), .Z(n208) );
  IV I_20 ( .A(TXELECIDLE), .Z(n209) );
  IV I_19 ( .A(n211), .Z(n210) );
  OR2 C240 ( .A(TXDATA[0]), .B(n212), .Z(n211) );
  OR2 C239 ( .A(n225), .B(n229), .Z(n212) );
  IV I_18 ( .A(n214), .Z(n213) );
  OR2 C225 ( .A(n224), .B(n228), .Z(n214) );
  IV I_17 ( .A(n216), .Z(n215) );
  OR2 C210 ( .A(n224), .B(n217), .Z(n216) );
  OR2 C209 ( .A(n225), .B(n218), .Z(n217) );
  OR2 C208 ( .A(TXDATA[2]), .B(n230), .Z(n218) );
  IV I_16 ( .A(n220), .Z(n219) );
  OR2 C195 ( .A(n224), .B(n221), .Z(n220) );
  OR2 C194 ( .A(n225), .B(n222), .Z(n221) );
  OR2 C193 ( .A(n282), .B(n223), .Z(n222) );
  OR2 C192 ( .A(TXDATA[3]), .B(n231), .Z(n223) );
  IV I_15 ( .A(TXDATA[0]), .Z(n224) );
  IV I_14 ( .A(TXDATA[1]), .Z(n225) );
  IV I_13 ( .A(n227), .Z(n226) );
  OR2 C180 ( .A(TXDATA[0]), .B(n228), .Z(n227) );
  OR2 C179 ( .A(TXDATA[1]), .B(n229), .Z(n228) );
  OR2 C178 ( .A(n282), .B(n230), .Z(n229) );
  OR2 C177 ( .A(n283), .B(n231), .Z(n230) );
  OR2 C176 ( .A(n284), .B(n232), .Z(n231) );
  OR2 C175 ( .A(n273), .B(n240), .Z(n232) );
  IV I_12 ( .A(n234), .Z(n233) );
  OR2 C166 ( .A(TXDATA[0]), .B(n235), .Z(n234) );
  OR2 C165 ( .A(TXDATA[1]), .B(n236), .Z(n235) );
  OR2 C164 ( .A(n282), .B(n237), .Z(n236) );
  OR2 C163 ( .A(n283), .B(n238), .Z(n237) );
  OR2 C162 ( .A(n284), .B(n239), .Z(n238) );
  OR2 C161 ( .A(TXDATA[5]), .B(n240), .Z(n239) );
  OR2 C160 ( .A(n265), .B(n256), .Z(n240) );
  IV I_11 ( .A(n242), .Z(n241) );
  OR2 C153 ( .A(TXDATA[0]), .B(n243), .Z(n242) );
  OR2 C152 ( .A(TXDATA[1]), .B(n244), .Z(n243) );
  OR2 C151 ( .A(n282), .B(n245), .Z(n244) );
  OR2 C150 ( .A(n283), .B(n246), .Z(n245) );
  OR2 C149 ( .A(n284), .B(n247), .Z(n246) );
  OR2 C148 ( .A(n273), .B(n255), .Z(n247) );
  IV I_10 ( .A(n249), .Z(n248) );
  OR2 C140 ( .A(TXDATA[0]), .B(n250), .Z(n249) );
  OR2 C139 ( .A(TXDATA[1]), .B(n251), .Z(n250) );
  OR2 C138 ( .A(n282), .B(n252), .Z(n251) );
  OR2 C137 ( .A(n283), .B(n253), .Z(n252) );
  OR2 C136 ( .A(n284), .B(n254), .Z(n253) );
  OR2 C135 ( .A(TXDATA[5]), .B(n255), .Z(n254) );
  OR2 C134 ( .A(TXDATA[6]), .B(n256), .Z(n255) );
  IV I_9 ( .A(TXDATA[7]), .Z(n256) );
  IV I_8 ( .A(n258), .Z(n257) );
  OR2 C128 ( .A(TXDATA[0]), .B(n259), .Z(n258) );
  OR2 C127 ( .A(TXDATA[1]), .B(n260), .Z(n259) );
  OR2 C126 ( .A(n282), .B(n261), .Z(n260) );
  OR2 C125 ( .A(n283), .B(n262), .Z(n261) );
  OR2 C124 ( .A(n284), .B(n263), .Z(n262) );
  OR2 C123 ( .A(TXDATA[5]), .B(n264), .Z(n263) );
  OR2 C122 ( .A(n265), .B(TXDATA[7]), .Z(n264) );
  IV I_7 ( .A(TXDATA[6]), .Z(n265) );
  IV I_6 ( .A(n267), .Z(n266) );
  OR2 C116 ( .A(TXDATA[0]), .B(n268), .Z(n267) );
  OR2 C115 ( .A(TXDATA[1]), .B(n269), .Z(n268) );
  OR2 C114 ( .A(n282), .B(n270), .Z(n269) );
  OR2 C113 ( .A(n283), .B(n271), .Z(n270) );
  OR2 C112 ( .A(n284), .B(n272), .Z(n271) );
  OR2 C111 ( .A(n273), .B(n281), .Z(n272) );
  IV I_5 ( .A(TXDATA[5]), .Z(n273) );
  IV I_4 ( .A(n275), .Z(n274) );
  OR2 C104 ( .A(TXDATA[0]), .B(n276), .Z(n275) );
  OR2 C103 ( .A(TXDATA[1]), .B(n277), .Z(n276) );
  OR2 C102 ( .A(n282), .B(n278), .Z(n277) );
  OR2 C101 ( .A(n283), .B(n279), .Z(n278) );
  OR2 C100 ( .A(n284), .B(n280), .Z(n279) );
  OR2 C99 ( .A(TXDATA[5]), .B(n281), .Z(n280) );
  OR2 C98 ( .A(TXDATA[6]), .B(TXDATA[7]), .Z(n281) );
  IV I_3 ( .A(TXDATA[2]), .Z(n282) );
  IV I_2 ( .A(TXDATA[3]), .Z(n283) );
  IV I_1 ( .A(TXDATA[4]), .Z(n284) );
  IV I_0 ( .A(TXDATAK), .Z(n285) );
  FD1 InputDataK_P0_reg ( .D(n511), .CP(PCLK250), .Q(n312) );
  FD1 InputCompliance_P0_reg ( .D(n510), .CP(PCLK250), .Q(n311) );
  FD1 InputData_P0_reg_7_ ( .D(n509), .CP(PCLK250), .Q(n320) );
  FD1 InputData_P0_reg_6_ ( .D(n508), .CP(PCLK250), .Q(n319) );
  FD1 InputData_P0_reg_5_ ( .D(n507), .CP(PCLK250), .Q(n318) );
  FD1 InputData_P0_reg_4_ ( .D(n506), .CP(PCLK250), .Q(n317) );
  FD1 InputData_P0_reg_3_ ( .D(n505), .CP(PCLK250), .Q(n316) );
  FD1 InputData_P0_reg_2_ ( .D(n504), .CP(PCLK250), .Q(n315) );
  FD1 InputData_P0_reg_1_ ( .D(n503), .CP(PCLK250), .Q(n314) );
  FD1 InputData_P0_reg_0_ ( .D(n502), .CP(PCLK250), .Q(n313) );
  FD1 InputDataEnable_P0_reg ( .D(U7_Z_0), .CP(PCLK250), .Q(n310) );
  FD1 OutputElecIdle_P0_reg ( .D(U5_Z_0), .CP(PCLK250), .Q(HSS_TXELECIDLE) );
  FD1 DISPARITY_P0_reg ( .D(n5), .CP(PCLK250), .Q(n4) );
  FD1 OutputData_P0_reg_7_ ( .D(n501), .CP(PCLK250), .Q(HSS_TXD[7]) );
  FD1 OutputData_P0_reg_8_ ( .D(n500), .CP(PCLK250), .Q(HSS_TXD[8]) );
  FD1 OutputData_P0_reg_4_ ( .D(n499), .CP(PCLK250), .Q(HSS_TXD[4]) );
  FD1 OutputData_P0_reg_9_ ( .D(n498), .CP(PCLK250), .Q(HSS_TXD[9]) );
  FD1 OutputData_P0_reg_6_ ( .D(n497), .CP(PCLK250), .Q(HSS_TXD[6]) );
  FD1 OutputData_P0_reg_5_ ( .D(n496), .CP(PCLK250), .Q(HSS_TXD[5]) );
  FD1 OutputData_P0_reg_0_ ( .D(n495), .CP(PCLK250), .Q(HSS_TXD[0]) );
  FD1 OutputData_P0_reg_1_ ( .D(n494), .CP(PCLK250), .Q(HSS_TXD[1]) );
  FD1 OutputData_P0_reg_2_ ( .D(n493), .CP(PCLK250), .Q(HSS_TXD[2]) );
  FD1 OutputData_P0_reg_3_ ( .D(n492), .CP(PCLK250), .Q(HSS_TXD[3]) );
  AN2 U34 ( .A(RX_LoopbackData_P2[0]), .B(CNTL_Loopback_P0), .Z(n399) );
  AN2 U92 ( .A(U7_DATA2_0), .B(TXDATA[0]), .Z(n446) );
  AN2 U95 ( .A(TXDATA[1]), .B(U7_DATA2_0), .Z(n449) );
  AN2 U98 ( .A(TXDATA[2]), .B(U7_DATA2_0), .Z(n451) );
  AN2 U101 ( .A(TXDATA[3]), .B(U7_DATA2_0), .Z(n453) );
  AN2 U104 ( .A(TXDATA[4]), .B(U7_DATA2_0), .Z(n455) );
  AN2 U107 ( .A(TXDATA[5]), .B(U7_DATA2_0), .Z(n457) );
  AN2 U110 ( .A(TXDATA[6]), .B(U7_DATA2_0), .Z(n459) );
  AN2 U113 ( .A(TXDATA[7]), .B(U7_DATA2_0), .Z(n461) );
  AN2 U116 ( .A(TXCOMPLIANCE), .B(U7_DATA2_0), .Z(n463) );
  IV U119 ( .A(U7_DATA2_0), .Z(n448) );
  AN2 U120 ( .A(TXDATAK), .B(U7_DATA2_0), .Z(n465) );
  AN2 U187 ( .A(CNTL_RESETN_P0), .B(U7_DATA2_0), .Z(U7_Z_0) );
  IV U200 ( .A(n45), .Z(n549) );
  IV U201 ( .A(n48), .Z(n548) );
  IV U202 ( .A(n72), .Z(n547) );
  IV U203 ( .A(n85), .Z(n546) );
  IV U204 ( .A(n89), .Z(n545) );
  IV U205 ( .A(n93), .Z(n544) );
  IV U206 ( .A(n75), .Z(n542) );
  IV U207 ( .A(n98), .Z(n541) );
  IV U208 ( .A(n100), .Z(n540) );
  IV U209 ( .A(n102), .Z(n539) );
  IV U210 ( .A(n104), .Z(n538) );
  IV U211 ( .A(n106), .Z(n537) );
  IV U212 ( .A(n108), .Z(n536) );
  IV U213 ( .A(n111), .Z(n535) );
  IV U214 ( .A(n78), .Z(n533) );
  IV U215 ( .A(n113), .Z(n532) );
  IV U216 ( .A(n115), .Z(n531) );
  IV U217 ( .A(n118), .Z(n530) );
  IV U218 ( .A(n122), .Z(n529) );
  IV U219 ( .A(n126), .Z(n528) );
  IV U220 ( .A(n130), .Z(n527) );
  IV U221 ( .A(n132), .Z(n526) );
  IV U222 ( .A(n30), .Z(n525) );
  IV U223 ( .A(n39), .Z(n522) );
  IV U224 ( .A(n54), .Z(n521) );
  IV U225 ( .A(n66), .Z(n520) );
  IV U226 ( .A(n70), .Z(n519) );
  IV U227 ( .A(n57), .Z(n517) );
  IV U228 ( .A(n311), .Z(n516) );
  IV U229 ( .A(n50), .Z(n513) );
  IV U230 ( .A(n24), .Z(n512) );
  OR2 U231 ( .A(n557), .B(n465), .Z(n511) );
  AN2 U232 ( .A(n448), .B(n312), .Z(n557) );
  OR2 U233 ( .A(n558), .B(n463), .Z(n510) );
  AN2 U234 ( .A(n448), .B(n311), .Z(n558) );
  OR2 U235 ( .A(n559), .B(n461), .Z(n509) );
  AN2 U236 ( .A(n448), .B(n320), .Z(n559) );
  OR2 U237 ( .A(n560), .B(n459), .Z(n508) );
  AN2 U238 ( .A(n448), .B(n319), .Z(n560) );
  OR2 U239 ( .A(n561), .B(n457), .Z(n507) );
  AN2 U240 ( .A(n448), .B(n318), .Z(n561) );
  OR2 U241 ( .A(n562), .B(n455), .Z(n506) );
  AN2 U242 ( .A(n448), .B(n317), .Z(n562) );
  OR2 U243 ( .A(n563), .B(n453), .Z(n505) );
  AN2 U244 ( .A(n448), .B(n316), .Z(n563) );
  OR2 U245 ( .A(n564), .B(n451), .Z(n504) );
  AN2 U246 ( .A(n448), .B(n315), .Z(n564) );
  OR2 U247 ( .A(n565), .B(n449), .Z(n503) );
  AN2 U248 ( .A(n448), .B(n314), .Z(n565) );
  OR2 U249 ( .A(n566), .B(n446), .Z(n502) );
  AN2 U250 ( .A(n448), .B(n313), .Z(n566) );
  OR2 U251 ( .A(n567), .B(n568), .Z(n501) );
  OR2 U252 ( .A(n569), .B(n570), .Z(n568) );
  AN2 U253 ( .A(HSS_TXD[7]), .B(n571), .Z(n570) );
  AN2 U254 ( .A(RX_LoopbackData_P2[7]), .B(n572), .Z(n569) );
  OR2 U255 ( .A(n573), .B(n574), .Z(n567) );
  AN2 U256 ( .A(n575), .B(n26), .Z(n574) );
  AN2 U257 ( .A(n576), .B(n577), .Z(n573) );
  IV U258 ( .A(n26), .Z(n577) );
  OR2 U259 ( .A(n578), .B(n579), .Z(n500) );
  OR2 U260 ( .A(n580), .B(n581), .Z(n579) );
  AN2 U261 ( .A(HSS_TXD[8]), .B(n571), .Z(n581) );
  AN2 U262 ( .A(RX_LoopbackData_P2[8]), .B(n572), .Z(n580) );
  OR2 U263 ( .A(n582), .B(n583), .Z(n578) );
  AN2 U264 ( .A(n575), .B(n320), .Z(n583) );
  AN2 U265 ( .A(n576), .B(n518), .Z(n582) );
  IV U266 ( .A(n320), .Z(n518) );
  OR2 U267 ( .A(n584), .B(n585), .Z(n499) );
  OR2 U268 ( .A(n586), .B(n587), .Z(n585) );
  AN2 U269 ( .A(n588), .B(U4_DATA2_4), .Z(n587) );
  AN2 U270 ( .A(RX_LoopbackData_P2[4]), .B(n572), .Z(n586) );
  AN2 U271 ( .A(HSS_TXD[4]), .B(n571), .Z(n584) );
  OR2 U272 ( .A(n589), .B(n590), .Z(n498) );
  OR2 U273 ( .A(n591), .B(n592), .Z(n590) );
  AN2 U274 ( .A(HSS_TXD[9]), .B(n571), .Z(n592) );
  AN2 U275 ( .A(RX_LoopbackData_P2[9]), .B(n572), .Z(n591) );
  OR2 U276 ( .A(n593), .B(n594), .Z(n589) );
  AN2 U277 ( .A(n27), .B(n575), .Z(n594) );
  AN2 U278 ( .A(n576), .B(n595), .Z(n593) );
  IV U279 ( .A(n27), .Z(n595) );
  OR2 U280 ( .A(n596), .B(n597), .Z(n497) );
  OR2 U281 ( .A(n598), .B(n599), .Z(n597) );
  AN2 U282 ( .A(HSS_TXD[6]), .B(n571), .Z(n599) );
  AN2 U283 ( .A(RX_LoopbackData_P2[6]), .B(n572), .Z(n598) );
  OR2 U284 ( .A(n600), .B(n601), .Z(n596) );
  AN2 U285 ( .A(n25), .B(n575), .Z(n601) );
  AN2 U286 ( .A(n602), .B(n588), .Z(n575) );
  IV U287 ( .A(n33), .Z(n602) );
  AN2 U288 ( .A(n576), .B(n603), .Z(n600) );
  IV U289 ( .A(n25), .Z(n603) );
  AN2 U290 ( .A(n588), .B(n33), .Z(n576) );
  OR2 U291 ( .A(n604), .B(n605), .Z(n496) );
  OR2 U292 ( .A(n606), .B(n607), .Z(n605) );
  AN2 U293 ( .A(n588), .B(U4_DATA2_5), .Z(n607) );
  AN2 U294 ( .A(RX_LoopbackData_P2[5]), .B(n572), .Z(n606) );
  AN2 U295 ( .A(HSS_TXD[5]), .B(n571), .Z(n604) );
  OR2 U296 ( .A(n608), .B(n609), .Z(n495) );
  AN2 U297 ( .A(n310), .B(n610), .Z(n609) );
  OR2 U298 ( .A(n611), .B(n399), .Z(n610) );
  AN2 U299 ( .A(n208), .B(n612), .Z(n611) );
  OR2 U300 ( .A(n34), .B(n613), .Z(n612) );
  OR2 U301 ( .A(n614), .B(n615), .Z(n613) );
  AN2 U302 ( .A(n313), .B(n616), .Z(n615) );
  AN2 U303 ( .A(n32), .B(n552), .Z(n614) );
  AN2 U304 ( .A(HSS_TXD[0]), .B(n571), .Z(n608) );
  OR2 U305 ( .A(n617), .B(n618), .Z(n494) );
  OR2 U306 ( .A(n619), .B(n620), .Z(n618) );
  AN2 U307 ( .A(HSS_TXD[1]), .B(n571), .Z(n620) );
  AN2 U308 ( .A(RX_LoopbackData_P2[1]), .B(n572), .Z(n619) );
  OR2 U309 ( .A(n621), .B(n622), .Z(n617) );
  AN2 U310 ( .A(n623), .B(n[6]), .Z(n622) );
  AN2 U311 ( .A(n624), .B(n625), .Z(n621) );
  IV U312 ( .A(n[6]), .Z(n625) );
  OR2 U313 ( .A(n626), .B(n627), .Z(n493) );
  OR2 U314 ( .A(n628), .B(n629), .Z(n627) );
  AN2 U315 ( .A(HSS_TXD[2]), .B(n571), .Z(n629) );
  AN2 U316 ( .A(RX_LoopbackData_P2[2]), .B(n572), .Z(n628) );
  OR2 U317 ( .A(n630), .B(n631), .Z(n626) );
  AN2 U318 ( .A(n[7]), .B(n623), .Z(n631) );
  AN2 U319 ( .A(n624), .B(n632), .Z(n630) );
  IV U320 ( .A(n[7]), .Z(n632) );
  OR2 U321 ( .A(n633), .B(n634), .Z(n492) );
  OR2 U322 ( .A(n635), .B(n636), .Z(n634) );
  AN2 U323 ( .A(HSS_TXD[3]), .B(n571), .Z(n636) );
  AN2 U324 ( .A(RX_LoopbackData_P2[3]), .B(n572), .Z(n635) );
  AN2 U325 ( .A(n310), .B(CNTL_Loopback_P0), .Z(n572) );
  OR2 U326 ( .A(n637), .B(n638), .Z(n633) );
  AN2 U327 ( .A(n[8]), .B(n623), .Z(n638) );
  AN2 U328 ( .A(n616), .B(n588), .Z(n623) );
  AN2 U329 ( .A(n624), .B(n639), .Z(n637) );
  IV U330 ( .A(n[8]), .Z(n639) );
  AN2 U331 ( .A(n588), .B(n32), .Z(n624) );
  AN2 U332 ( .A(n208), .B(n640), .Z(n588) );
  IV U333 ( .A(n641), .Z(n640) );
  OR2 U334 ( .A(n34), .B(n571), .Z(n641) );
  OR2 U335 ( .A(n642), .B(n643), .Z(n178) );
  IV U336 ( .A(n644), .Z(n643) );
  OR2 U337 ( .A(n514), .B(n177), .Z(n644) );
  AN2 U338 ( .A(n177), .B(n514), .Z(n642) );
  IV U339 ( .A(n23), .Z(n514) );
  OR2 U340 ( .A(n645), .B(n646), .Z(n23) );
  AN2 U341 ( .A(n175), .B(n515), .Z(n646) );
  IV U342 ( .A(n647), .Z(n645) );
  OR2 U343 ( .A(n515), .B(n175), .Z(n647) );
  IV U344 ( .A(n31), .Z(n515) );
  OR2 U345 ( .A(n648), .B(n649), .Z(n171) );
  AN2 U346 ( .A(n318), .B(n523), .Z(n649) );
  IV U347 ( .A(n319), .Z(n523) );
  AN2 U348 ( .A(n319), .B(n524), .Z(n648) );
  IV U349 ( .A(n318), .Z(n524) );
  OR2 U350 ( .A(n650), .B(n651), .Z(n143) );
  AN2 U351 ( .A(n315), .B(n543), .Z(n651) );
  IV U352 ( .A(n316), .Z(n543) );
  AN2 U353 ( .A(n316), .B(n550), .Z(n650) );
  IV U354 ( .A(n315), .Z(n550) );
  OR2 U355 ( .A(n652), .B(n653), .Z(n142) );
  AN2 U356 ( .A(n313), .B(n551), .Z(n653) );
  IV U357 ( .A(n314), .Z(n551) );
  AN2 U358 ( .A(n314), .B(n552), .Z(n652) );
  IV U359 ( .A(n313), .Z(n552) );
  OR2 U360 ( .A(n654), .B(n655), .Z(n140) );
  IV U361 ( .A(n656), .Z(n655) );
  OR2 U362 ( .A(n534), .B(n43), .Z(n656) );
  AN2 U363 ( .A(n43), .B(n534), .Z(n654) );
  AN2 U364 ( .A(n657), .B(n658), .Z(n137) );
  IV U365 ( .A(n659), .Z(n658) );
  AN2 U366 ( .A(n534), .B(n81), .Z(n659) );
  OR2 U367 ( .A(n81), .B(n534), .Z(n657) );
  IV U368 ( .A(n317), .Z(n534) );
  OR2 U369 ( .A(n660), .B(n207), .Z(U5_Z_0) );
  AN2 U370 ( .A(CNTL_RESETN_P0), .B(n571), .Z(n660) );
  IV U371 ( .A(n310), .Z(n571) );
  OR2 U372 ( .A(n661), .B(n662), .Z(U4_DATA2_5) );
  AN2 U373 ( .A(n[10]), .B(n616), .Z(n662) );
  IV U374 ( .A(n663), .Z(n661) );
  OR2 U375 ( .A(n616), .B(n[10]), .Z(n663) );
  OR2 U376 ( .A(n664), .B(n665), .Z(U4_DATA2_4) );
  IV U377 ( .A(n666), .Z(n665) );
  OR2 U378 ( .A(n616), .B(n[9]), .Z(n666) );
  AN2 U379 ( .A(n[9]), .B(n616), .Z(n664) );
  IV U380 ( .A(n32), .Z(n616) );
endmodule

