
module XFIPCS_TX_PCS ( pma_tx_clk, reset_to_pma_tx, reset_to_xgmii_tx, 
        enable_alternate_refresh, ALTERNATE_ENCODE, loopback_xgmii, txc_xfi, 
        txd_xfi, tx_fifo_pop_pre, test_pat_seed_a, test_pat_seed_b, 
        tx_prbs_pat_en, tx_test_pat_en, test_pat_sel, data_pat_sel, 
        scr_bypass_enable, tx_data_out, tx_fifo_pop_2, tx_mode, t_type_li, 
        TXxQUIET, TXxREFRESH, assertion_shengyushen );
  input [7:0] txc_xfi;
  input [63:0] txd_xfi;
  input [57:0] test_pat_seed_a;
  input [57:0] test_pat_seed_b;
  output [65:0] tx_data_out;
  output [1:0] tx_mode;
  input pma_tx_clk, reset_to_pma_tx, reset_to_xgmii_tx,
         enable_alternate_refresh, ALTERNATE_ENCODE, loopback_xgmii,
         tx_fifo_pop_pre, tx_prbs_pat_en, tx_test_pat_en, test_pat_sel,
         data_pat_sel, scr_bypass_enable;
  output tx_fifo_pop_2, t_type_li, TXxQUIET, TXxREFRESH, assertion_shengyushen;
  wire   n32, n35, n38, n41, n44, n97, n98, n99, n110, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n143, n159, n175, n191, n207, n223,
         n239, n255, n257, n259, n261, n263, n265, n267, n269, n271, n273,
         n275, n277, n279, n281, n283, n285, n287, n289, n291, n293, n295,
         n297, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n324, n325, n326, n327, n328, n331, n334, n335,
         n336, n338, n339, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n749, n750, n816, n817, n940, n1115, n1148, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1459, n1460, n1461, n1462, n1465,
         n1466, n1467, n1468, n1471, n1472, n1473, n1474, n1477, n1478, n1479,
         n1480, n1483, n1484, n1485, n1486, n1489, n1490, n1491, n1492, n1495,
         n1496, n1497, n1498, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1509, n1510, n1511, n1512, n1514, n1515, n1516, n1517, n1518, n1519,
         n1521, n1522, n1523, n1524, n1525, n1526, n1528, n1529, n1530, n1531,
         n1532, n1533, n1535, n1536, n1537, n1538, n1539, n1540, n1542, n1543,
         n1544, n1545, n1546, n1547, n1549, n1550, n1551, n1552, n1553, n1554,
         n1556, n1557, n1558, n1559, n1560, n1561, n1563, n1564, n1565, n1566,
         n1567, n1568, n1570, n1571, n1572, n1573, n1574, n1575, n1577, n1578,
         n1579, n1580, n1581, n1582, n1584, n1585, n1586, n1587, n1588, n1589,
         n1591, n1592, n1593, n1594, n1595, n1596, n1598, n1599, n1600, n1601,
         n1602, n1603, n1605, n1606, n1607, n1608, n1609, n1610, n1612, n1613,
         n1614, n1615, n1616, n1617, n1619, n1620, n1621, n1622, n1623, n1624,
         n1626, n1627, n1628, n1629, n1630, n1632, n1633, n1634, n1635, n1636,
         n1638, n1639, n1640, n1641, n1642, n1644, n1645, n1646, n1647, n1648,
         n1650, n1651, n1652, n1653, n1654, n1656, n1657, n1658, n1659, n1660,
         n1662, n1663, n1664, n1665, n1666, n1668, n1669, n1670, n1671, n1672,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1778, n1779, n1780, n1781, n1782, n1783, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1793, n1794, n1795, n1796, n1797, n1798,
         n1800, n1803, n1806, n1809, n1812, n1815, n1818, n1821, n1824, n1825,
         n1827, n1828, n1830, n1831, n1833, n1834, n1836, n1837, n1839, n1840,
         n1842, n1843, n1845, n1846, n1848, n1849, n1850, n1852, n1853, n1854,
         n1855, n1856, n1857, n1859, n1860, n1861, n1863, n1864, n1865, n1866,
         n1867, n1868, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1905, n1906, n1907, n1909, n1910, n1914,
         n1918, n1919, n1924, n1926, n1927, n1929, n1930, n1932, n1934, n1935,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2516, n2517, n2533, n2534, n2536, n2537, n2540, n2541, n2544,
         n2545, n2548, n2549, n2551, n2552, n2555, n2556, n2559, n2560, n2563,
         n2564, n2566, n2567, n2569, n2570, n2572, n2573, n2575, n2576, n2578,
         n2579, n2581, n2582, n2584, n2585, n2587, n2593, n2664, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2747, n2749, n2753,
         n2756, n2757, n2760, n2762, n2770, n2771, n2774, n2775, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2861, n2862,
         n2863, n2864, n2867, n2868, n2871, n2872, n2875, n2876, n2879, n2880,
         n2884, n2892, n2900, n2915, n2923, n2937, n2946, n2947, n2948, n2951,
         n2952, n2953, n2956, n2957, n2958, n2960, n2961, n2963, n2964, n2966,
         n2967, n2968, n2972, n2974, n2975, n2977, n2979, n2985, n2987, n2988,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3179, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3267, n3268, n3271, n3272, n3273,
         n3279, n3281, n3284, n3286, n3288, n3290, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3431, n3432, n3433, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3476, n3477, n3478,
         n3479, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3497, n3498, n3499, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3519, n3520, n3521, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4170, n4172, n4173, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4369, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4475, n4476, n4477,
         n4479, n4480, n4614, U3_U1_Z_1, U3_U1_Z_2, U3_U1_Z_3, U3_U1_Z_4,
         U3_U1_Z_5, U3_U1_Z_6, U3_U1_Z_7, U3_U1_Z_8, U3_U1_Z_9, U3_U1_Z_10,
         U3_U1_Z_11, U3_U1_Z_12, U3_U1_Z_13, U3_U1_Z_14, U3_U1_Z_15,
         U3_U1_DATA3_0, U3_U1_DATA3_1, U3_U1_DATA3_2, U3_U1_DATA3_3,
         U3_U1_DATA3_4, U3_U1_DATA3_5, U3_U1_DATA3_6, U3_U1_DATA3_7,
         U3_U1_DATA3_8, U3_U1_DATA3_9, U3_U1_DATA3_10, U3_U1_DATA1_0,
         U3_U1_DATA1_1, U3_U1_DATA1_2, U3_U1_DATA1_3, U3_U1_DATA1_4,
         U3_U1_DATA1_5, U3_U1_DATA1_6, U3_U1_DATA1_7, U3_U1_DATA1_8,
         U3_U1_DATA1_9, U3_U1_DATA1_10, U3_U1_DATA1_11, U3_U1_DATA1_12,
         U3_U1_DATA1_13, U3_U1_DATA1_14, U3_U1_DATA1_15, U162_Z_0, U162_Z_1,
         U162_Z_2, U162_Z_3, U162_Z_4, U162_Z_5, U162_Z_6, U162_Z_7, U162_Z_8,
         U162_Z_9, U162_Z_10, U162_Z_11, U162_Z_12, U162_Z_13, U162_Z_14,
         U162_Z_15, U162_Z_16, U162_Z_17, U162_Z_18, U162_Z_19, U162_Z_20,
         U162_Z_21, U162_Z_22, U162_Z_23, U162_Z_24, U162_Z_25, U162_Z_26,
         U162_Z_27, U162_Z_28, U162_Z_29, U162_Z_30, U162_Z_31, U162_Z_32,
         U162_Z_33, U162_Z_34, U162_Z_35, U162_Z_36, U162_Z_37, U162_Z_38,
         U162_Z_39, U162_Z_40, U162_Z_41, U162_Z_42, U162_Z_43, U162_Z_44,
         U162_Z_45, U162_Z_46, U162_Z_47, U162_Z_48, U162_Z_49, U162_Z_50,
         U162_Z_51, U162_Z_52, U162_Z_53, U162_Z_54, U162_Z_55, U162_Z_56,
         U162_Z_57, U162_Z_58, U162_Z_59, U162_Z_60, U162_Z_61, U162_Z_62,
         U162_Z_63, U162_DATA3_0, U162_DATA3_1, U162_DATA3_2, U162_DATA3_3,
         U162_DATA3_4, U162_DATA3_5, U162_DATA3_6, U162_DATA3_7, U162_DATA3_8,
         U162_DATA3_9, U162_DATA3_10, U162_DATA3_11, U162_DATA3_12,
         U162_DATA3_13, U162_DATA3_14, U162_DATA3_15, U162_DATA3_16,
         U162_DATA3_17, U162_DATA3_18, U162_DATA3_19, U162_DATA3_20,
         U162_DATA3_21, U162_DATA3_22, U162_DATA3_23, U162_DATA3_24,
         U162_DATA3_25, U162_DATA3_26, U162_DATA3_27, U162_DATA3_28,
         U162_DATA3_29, U162_DATA3_30, U162_DATA3_31, U162_DATA3_32,
         U162_DATA3_33, U162_DATA3_34, U162_DATA3_35, U162_DATA3_36,
         U162_DATA3_37, U162_DATA3_38, U162_DATA3_39, U162_DATA3_40,
         U162_DATA3_41, U162_DATA3_42, U162_DATA3_43, U162_DATA3_44,
         U162_DATA3_45, U162_DATA3_46, U162_DATA3_47, U162_DATA3_48,
         U162_DATA3_49, U162_DATA3_50, U162_DATA3_51, U162_DATA3_52,
         U162_DATA3_53, U162_DATA3_54, U162_DATA3_55, U162_DATA3_56,
         U162_DATA3_57, U162_DATA3_58, U162_DATA3_59, U162_DATA3_60,
         U162_DATA3_61, U162_DATA3_62, U162_DATA3_63, U161_Z_0, U161_Z_1,
         U161_Z_2, U161_Z_3, U161_Z_4, U161_Z_5, U161_Z_6, U161_Z_7,
         U161_CONTROL3, U161_CONTROL2, U161_DATA3_0, U161_DATA3_1,
         U161_DATA3_2, U161_DATA3_3, U161_DATA3_4, U161_DATA3_5, U161_DATA3_6,
         U161_DATA3_7, U160_Z_0, U160_Z_1, U160_Z_2, U160_Z_3, U160_DATA2_0,
         U160_DATA2_1, U160_DATA2_2, U160_DATA2_3, U159_Z_0, U159_Z_1,
         U159_Z_2, U159_Z_3, U159_Z_4, U159_Z_5, U159_Z_6, U159_Z_7, U158_Z_0,
         U158_Z_1, U158_Z_3, U158_Z_5, U158_Z_6, U158_Z_8, U158_Z_9, U158_Z_11,
         U158_Z_13, U158_Z_14, U157_Z_0, U157_Z_1, U157_Z_2, U157_Z_3,
         U157_Z_4, U157_Z_5, U157_CONTROL2, U156_Z_0, U156_Z_1, U156_Z_2,
         U156_Z_3, U156_Z_4, U156_Z_5, U156_Z_6, U156_Z_7, U156_Z_8, U156_Z_9,
         U156_Z_10, U156_Z_11, U156_Z_12, U156_Z_13, U156_Z_14, U156_Z_15,
         U156_Z_16, U156_Z_17, U156_Z_18, U156_Z_19, U156_Z_20, U156_Z_21,
         U156_Z_22, U156_Z_23, U156_Z_24, U156_Z_25, U156_Z_26, U156_Z_27,
         U156_Z_28, U156_Z_29, U156_Z_30, U156_Z_31, U156_Z_32, U156_Z_33,
         U155_Z_0, U155_Z_1, U154_Z_0, U154_Z_1, U154_Z_2, U154_Z_3, U154_Z_4,
         U154_Z_5, U153_DATA2_0, U152_DATA3_0, U151_DATA3_0, U150_DATA3_0,
         U149_DATA2_0, U148_DATA3_0, U141_CONTROL2, U140_CONTROL2,
         U124_CONTROL2, U122_CONTROL2, U119_Z_0, U119_Z_1, U119_Z_2, U119_Z_3,
         U118_Z_0, U118_Z_1, U117_Z_0, U117_Z_1, U117_Z_2, U117_Z_3, U117_Z_4,
         U117_Z_5, U117_Z_6, U117_Z_7, U117_Z_8, U117_Z_9, U117_Z_10,
         U117_Z_11, U117_Z_12, U117_Z_13, U117_Z_14, U117_Z_15, U114_DATA2_0,
         U113_DATA3_0, U112_DATA3_0, U111_DATA3_0, U107_DATA1_0, U76_DATA4_0,
         U76_DATA3_0, U73_DATA6_0, U73_DATA5_0, U72_DATA3_0, U72_DATA2_0,
         U71_DATA3_0, U69_DATA4_0, U69_DATA2_0, U67_Z_0, U67_Z_1, U67_Z_2,
         U67_Z_3, U66_Z_0, U66_Z_1, U65_Z_0, U64_Z_0, U63_Z_0, U61_DATA2_1,
         U61_DATA2_2, U61_DATA2_8, U61_DATA2_9, U61_DATA2_15, U61_DATA2_16,
         U61_DATA2_22, U61_DATA2_23, U59_DATA1_0, U59_DATA1_1, U57_DATA1_0,
         U57_DATA1_1, U55_DATA1_1, U54_DATA1_0, U52_DATA1_1, U52_DATA1_2,
         U40_DATA2_0, U40_DATA2_1, U40_DATA2_2, U40_DATA2_3, U40_DATA2_4,
         U40_DATA2_5, U40_DATA2_6, U40_DATA2_7, U37_DATA6_0, U37_DATA6_1,
         U37_DATA6_2, U37_DATA6_3, U37_DATA6_4, U37_DATA6_5, U37_DATA6_6,
         U37_DATA6_7, U37_DATA6_8, U37_DATA6_9, U37_DATA6_10, U37_DATA6_11,
         U37_DATA6_12, U37_DATA6_13, U37_DATA6_14, U37_DATA6_15, U37_DATA6_16,
         U37_DATA6_17, U37_DATA6_18, U37_DATA6_19, U37_DATA6_20, U37_DATA6_21,
         U37_DATA6_22, U37_DATA6_23, U37_DATA6_24, U37_DATA6_25, U37_DATA6_26,
         U37_DATA6_27, U37_DATA6_28, U37_DATA6_29, U37_DATA6_30, U37_DATA6_31,
         U37_DATA6_32, U37_DATA6_33, U37_DATA6_34, U37_DATA6_35, U37_DATA6_36,
         U37_DATA6_37, U37_DATA6_38, U37_DATA6_39, U37_DATA6_40, U37_DATA6_41,
         U37_DATA6_42, U37_DATA6_43, U37_DATA6_44, U37_DATA6_45, U37_DATA6_46,
         U37_DATA6_47, U37_DATA6_48, U37_DATA6_49, U37_DATA6_50, U37_DATA6_51,
         U37_DATA6_52, U37_DATA6_53, U37_DATA6_54, U37_DATA6_55, U37_DATA6_56,
         U37_DATA6_57, U37_DATA4_0, U37_DATA4_1, U37_DATA4_2, U37_DATA4_3,
         U37_DATA4_4, U37_DATA4_5, U37_DATA4_6, U37_DATA4_7, U37_DATA4_8,
         U37_DATA4_9, U37_DATA4_10, U37_DATA4_11, U37_DATA4_12, U37_DATA4_13,
         U37_DATA4_14, U37_DATA4_15, U37_DATA4_16, U37_DATA4_17, U37_DATA4_18,
         U37_DATA4_19, U37_DATA4_20, U37_DATA4_21, U37_DATA4_22, U37_DATA4_23,
         U37_DATA4_24, U37_DATA4_25, U37_DATA4_26, U37_DATA4_27, U37_DATA4_28,
         U37_DATA4_29, U37_DATA4_30, U37_DATA4_31, U37_DATA4_32, U37_DATA4_33,
         U37_DATA4_34, U37_DATA4_35, U37_DATA4_36, U37_DATA4_37, U37_DATA4_38,
         U37_DATA4_39, U37_DATA4_40, U37_DATA4_41, U37_DATA4_42, U37_DATA4_43,
         U37_DATA4_44, U37_DATA4_45, U37_DATA4_46, U37_DATA4_47, U37_DATA4_48,
         U37_DATA4_49, U37_DATA4_50, U37_DATA4_51, U37_DATA4_52, U37_DATA4_53,
         U37_DATA4_54, U37_DATA4_55, U37_DATA4_56, U37_DATA4_57, U37_DATA1_0,
         U37_DATA1_1, U37_DATA1_2, U37_DATA1_3, U37_DATA1_4, U37_DATA1_5,
         U37_DATA1_6, U37_DATA1_7, U37_DATA1_8, U37_DATA1_9, U37_DATA1_10,
         U37_DATA1_11, U37_DATA1_12, U37_DATA1_13, U37_DATA1_14, U37_DATA1_15,
         U37_DATA1_16, U37_DATA1_17, U37_DATA1_18, U37_DATA1_19, U37_DATA1_20,
         U37_DATA1_21, U37_DATA1_22, U37_DATA1_23, U37_DATA1_24, U37_DATA1_25,
         U37_DATA1_26, U37_DATA1_27, U37_DATA1_28, U37_DATA1_29, U37_DATA1_30,
         U37_DATA1_31, U37_DATA1_32, U37_DATA1_33, U37_DATA1_34, U37_DATA1_35,
         U37_DATA1_36, U37_DATA1_37, U37_DATA1_38, U37_DATA1_39, U37_DATA1_40,
         U37_DATA1_41, U37_DATA1_42, U37_DATA1_43, U37_DATA1_44, U37_DATA1_45,
         U37_DATA1_46, U37_DATA1_47, U37_DATA1_48, U37_DATA1_49, U37_DATA1_50,
         U37_DATA1_51, U37_DATA1_52, U37_DATA1_53, U37_DATA1_54, U37_DATA1_55,
         U37_DATA1_56, U37_DATA1_57, U35_Z_0, U35_Z_1, U35_Z_2, U35_Z_3,
         U35_Z_4, U35_Z_5, U35_Z_6, U35_Z_7, U35_Z_8, U35_Z_9, U35_Z_10,
         U35_Z_11, U35_Z_12, U35_Z_13, U35_Z_14, U35_Z_15, U35_Z_16, U35_Z_17,
         U35_Z_18, U35_Z_19, U35_Z_20, U35_Z_21, U35_Z_22, U35_Z_23, U35_Z_24,
         U35_Z_25, U35_Z_26, U35_Z_27, U35_Z_28, U35_Z_29, U35_Z_30, U35_Z_31,
         U35_Z_32, U35_Z_33, U35_Z_34, U35_Z_35, U35_Z_36, U35_Z_37, U35_Z_38,
         U35_Z_39, U35_Z_40, U35_Z_41, U35_Z_42, U35_Z_43, U35_Z_44, U35_Z_45,
         U35_Z_46, U35_Z_47, U35_Z_48, U35_Z_49, U35_Z_50, U35_Z_51, U35_Z_52,
         U35_Z_53, U35_Z_54, U35_Z_55, U35_Z_56, U35_Z_57, U34_Z_0, U34_Z_1,
         U34_Z_2, U34_Z_3, U34_Z_4, U34_Z_5, U34_Z_6, U34_Z_7, U34_Z_8, U8_Z_0,
         U8_Z_1, U8_Z_2, U8_Z_3, U8_Z_4, U8_Z_5, U8_Z_6, U8_Z_7, U8_Z_8,
         U8_Z_9, U8_Z_10, U7_Z_0, U7_Z_1, U7_Z_2, U7_Z_3, U7_Z_4, U7_Z_5,
         U7_Z_6, U7_Z_7, U7_Z_8, U7_Z_9, U7_Z_10, U7_Z_11, U7_Z_12, U7_Z_13,
         U7_Z_14, U7_Z_15, U7_Z_16, U7_Z_17, U7_Z_18, U7_Z_19, U6_Z_0, U6_Z_1,
         U6_Z_2, U6_Z_3, U6_Z_4, U6_Z_5, U6_Z_6, U6_Z_7, U6_Z_8, U6_Z_9,
         U6_Z_10, U6_Z_11, U5_Z_0, U5_Z_1, U5_Z_2, U5_Z_3, U5_Z_4, U5_Z_5,
         U5_Z_6, U5_Z_7, U5_Z_8, U4_DATA1_0, U4_DATA1_1, U4_DATA1_2,
         U4_DATA1_3, U4_DATA1_4, U4_DATA1_5, U4_DATA1_6, U4_DATA1_7,
         U4_DATA1_8, sub_128_aco_B_0_, sub_128_aco_A_0_, sub_128_aco_A_1_,
         sub_128_aco_A_2_, sub_128_aco_A_3_, sub_128_aco_A_4_,
         sub_128_aco_A_5_, sub_128_aco_A_6_, sub_128_aco_A_7_,
         sub_128_aco_A_8_, sub_127_aco_B_0_, sub_127_aco_A_0_,
         sub_127_aco_A_1_, sub_127_aco_A_2_, sub_127_aco_A_3_,
         sub_127_aco_A_4_, sub_127_aco_A_5_, sub_127_aco_A_6_,
         sub_127_aco_A_7_, sub_127_aco_A_8_, sub_127_aco_A_9_,
         sub_127_aco_A_10_, sub_127_aco_A_11_, sub_125_aco_B_0_, r224_GTV2_1_,
         r224_GTV2_2_, r224_GTV2_3_, r224_GTV2_4_, r224_GTV2_5_, r224_GTV2_6_,
         r224_GTV2_7_, r224_GTV2_8_, r224_GTV2_9_, r224_GTV2_10_,
         r224_GTV2_11_, r224_GTV2_12_, r224_GTV2_13_, r224_GTV2_14_,
         r224_GTV2_15_, r224_GTV_2_, r224_GTV_3_, r224_GTV_4_, r224_GTV_5_,
         r224_GTV_6_, r224_GTV_7_, r224_GTV_8_, r224_GTV_9_, r224_GTV_10_,
         r224_GTV_11_, r224_GTV_12_, r224_GTV_13_, r224_GTV_14_, r224_GTV_15_,
         r224_GT, sub_126_aco_B_0_, sub_126_aco_A_0_, sub_126_aco_A_1_,
         sub_126_aco_A_2_, sub_126_aco_A_3_, sub_126_aco_A_4_,
         sub_126_aco_A_5_, sub_126_aco_A_6_, sub_126_aco_A_7_,
         sub_126_aco_A_8_, sub_126_aco_A_9_, sub_126_aco_A_10_,
         sub_126_aco_A_11_, sub_126_aco_A_12_, sub_126_aco_A_13_,
         sub_126_aco_A_14_, sub_126_aco_A_15_, sub_126_aco_A_16_,
         sub_126_aco_A_17_, sub_126_aco_A_18_, sub_126_aco_A_19_, n4894, n4898,
         n4899, n4900, n4903, n4909, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4921, n4924, n4925, n4926, n4927, n4928, n4929, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5236, n5245, n5246, n5247, n5248,
         n5249, n5254, n5257, n5259, n5261, n5263, n5264, n5268, n5269, n5270,
         n5274, n5275, n5276, n5277, n5279, n5281, n5282, n5284, n5285, n5288,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5453, n5454,
         n5455, n5457, n5458, n5459, n5462, n5467, n5469, n5470, n5471, n5474,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5517, n5518,
         n5519, n5520, n5521, n5525, n5526, n5527, n5538, n5559, n5572, n5582,
         n5627, n5628, n5684, n5685, n8179, n8180, n8182, n8183, n8184, n8186,
         n8188, n8190, n8192, n8194, n8196, n8199, n8200, n8202, n8203, n8205,
         n8206, n8207, n8209, n8211, n8213, n8215, n8218, n8219, n8220, n8223,
         n8224, n8226, n8227, n8228, n8230, n8232, n8234, n8236, n8239, n8240,
         n8242, n8243, n8245, n8246, n8247, n8249, n8251, n8253, n8255, n8257,
         n8260, n8261, n8263, n8264, n8266, n8267, n8268, n8270, n8272, n8274,
         n8276, n8278, n8281, n8282, n8284, n8285, n8287, n8288, n8289, n8291,
         n8293, n8295, n8298, n8299, n8300, n8303, n8304, n8306, n8307, n8309,
         n8310, n8311, n8313, n8315, n8317, n8319, n8322, n8323, n8325, n8326,
         n8328, n8329, n8331, n8332, n8334, n8335, n8337, n8338, n8340, n8341,
         n8343, n8344, n8346, n8347, n8349, n8350, n8352, n8353, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853;
  wire   [3181:3184] n;

  OR2 r224_UGTI1 ( .A(U3_U1_Z_15), .B(n5487), .Z(r224_GTV2_15_) );
  OR2 r224_UGTI2 ( .A(U3_U1_Z_15), .B(n5486), .Z(r224_GT) );
  OR2 r224_UGTI1_1 ( .A(U3_U1_Z_1), .B(n5515), .Z(r224_GTV2_1_) );
  OR2 r224_UGTI2_1 ( .A(U3_U1_Z_1), .B(n5514), .Z(r224_GTV_2_) );
  OR2 r224_UGTI1_2 ( .A(U3_U1_Z_2), .B(n5513), .Z(r224_GTV2_2_) );
  OR2 r224_UGTI2_2 ( .A(U3_U1_Z_2), .B(n5512), .Z(r224_GTV_3_) );
  OR2 r224_UGTI1_3 ( .A(U3_U1_Z_3), .B(n5511), .Z(r224_GTV2_3_) );
  OR2 r224_UGTI2_3 ( .A(U3_U1_Z_3), .B(n5510), .Z(r224_GTV_4_) );
  OR2 r224_UGTI1_4 ( .A(U3_U1_Z_4), .B(n5509), .Z(r224_GTV2_4_) );
  OR2 r224_UGTI2_4 ( .A(U3_U1_Z_4), .B(n5508), .Z(r224_GTV_5_) );
  OR2 r224_UGTI1_5 ( .A(U3_U1_Z_5), .B(n5507), .Z(r224_GTV2_5_) );
  OR2 r224_UGTI2_5 ( .A(U3_U1_Z_5), .B(n5506), .Z(r224_GTV_6_) );
  OR2 r224_UGTI1_6 ( .A(U3_U1_Z_6), .B(n5505), .Z(r224_GTV2_6_) );
  OR2 r224_UGTI2_6 ( .A(U3_U1_Z_6), .B(n5504), .Z(r224_GTV_7_) );
  OR2 r224_UGTI1_7 ( .A(U3_U1_Z_7), .B(n5503), .Z(r224_GTV2_7_) );
  OR2 r224_UGTI2_7 ( .A(U3_U1_Z_7), .B(n5502), .Z(r224_GTV_8_) );
  OR2 r224_UGTI1_8 ( .A(U3_U1_Z_8), .B(n5501), .Z(r224_GTV2_8_) );
  OR2 r224_UGTI2_8 ( .A(U3_U1_Z_8), .B(n5500), .Z(r224_GTV_9_) );
  OR2 r224_UGTI1_9 ( .A(U3_U1_Z_9), .B(n5499), .Z(r224_GTV2_9_) );
  OR2 r224_UGTI2_9 ( .A(U3_U1_Z_9), .B(n5498), .Z(r224_GTV_10_) );
  OR2 r224_UGTI1_10 ( .A(U3_U1_Z_10), .B(n5497), .Z(r224_GTV2_10_) );
  OR2 r224_UGTI2_10 ( .A(U3_U1_Z_10), .B(n5496), .Z(r224_GTV_11_) );
  OR2 r224_UGTI1_11 ( .A(U3_U1_Z_11), .B(n5495), .Z(r224_GTV2_11_) );
  OR2 r224_UGTI2_11 ( .A(U3_U1_Z_11), .B(n5494), .Z(r224_GTV_12_) );
  OR2 r224_UGTI1_12 ( .A(U3_U1_Z_12), .B(n5493), .Z(r224_GTV2_12_) );
  OR2 r224_UGTI2_12 ( .A(U3_U1_Z_12), .B(n5492), .Z(r224_GTV_13_) );
  OR2 r224_UGTI1_13 ( .A(U3_U1_Z_13), .B(n5491), .Z(r224_GTV2_13_) );
  OR2 r224_UGTI2_13 ( .A(U3_U1_Z_13), .B(n5490), .Z(r224_GTV_14_) );
  OR2 r224_UGTI1_14 ( .A(U3_U1_Z_14), .B(n5489), .Z(r224_GTV2_14_) );
  OR2 r224_UGTI2_14 ( .A(U3_U1_Z_14), .B(n5488), .Z(r224_GTV_15_) );
  OR2 C949 ( .A(n5261), .B(n324), .Z(n408) );
  OR2 C950 ( .A(n325), .B(n326), .Z(n409) );
  OR2 C951 ( .A(n327), .B(n328), .Z(n410) );
  OR2 C952 ( .A(n5270), .B(n5281), .Z(n411) );
  OR2 C9531 ( .A(n331), .B(n5284), .Z(n412) );
  OR2 C9541 ( .A(n5279), .B(n334), .Z(n413) );
  OR2 C9551 ( .A(n335), .B(n336), .Z(n414) );
  OR2 C9561 ( .A(n408), .B(n409), .Z(n415) );
  OR2 C9571 ( .A(n410), .B(n411), .Z(n416) );
  OR2 C9581 ( .A(n412), .B(n413), .Z(n417) );
  OR2 C9591 ( .A(n414), .B(n8644), .Z(n418) );
  OR2 C960 ( .A(n415), .B(n416), .Z(n419) );
  OR2 C961 ( .A(n417), .B(n418), .Z(n420) );
  OR2 C9651 ( .A(n5261), .B(n324), .Z(n424) );
  OR2 C9661 ( .A(n325), .B(n326), .Z(n425) );
  OR2 C9671 ( .A(n327), .B(n328), .Z(n426) );
  OR2 C9681 ( .A(n5270), .B(n5281), .Z(n427) );
  OR2 C9691 ( .A(n331), .B(n5284), .Z(n428) );
  OR2 C9701 ( .A(n5279), .B(n334), .Z(n429) );
  OR2 C971 ( .A(n335), .B(n5285), .Z(n430) );
  OR2 C972 ( .A(n424), .B(n425), .Z(n431) );
  OR2 C973 ( .A(n426), .B(n427), .Z(n432) );
  OR2 C974 ( .A(n428), .B(n429), .Z(n433) );
  OR2 C975 ( .A(n430), .B(n5288), .Z(n434) );
  OR2 C976 ( .A(n431), .B(n432), .Z(n435) );
  OR2 C9771 ( .A(n433), .B(n434), .Z(n436) );
  OR2 C9811 ( .A(n5261), .B(n324), .Z(n440) );
  OR2 C9821 ( .A(n325), .B(n326), .Z(n441) );
  OR2 C9831 ( .A(n327), .B(n328), .Z(n442) );
  OR2 C984 ( .A(n5270), .B(n5281), .Z(n443) );
  OR2 C985 ( .A(n331), .B(n5284), .Z(n444) );
  OR2 C986 ( .A(n5279), .B(n334), .Z(n445) );
  OR2 C987 ( .A(n5276), .B(n336), .Z(n446) );
  OR2 C9881 ( .A(n440), .B(n441), .Z(n447) );
  OR2 C9891 ( .A(n442), .B(n443), .Z(n448) );
  OR2 C9901 ( .A(n444), .B(n445), .Z(n449) );
  OR2 C9911 ( .A(n446), .B(n5288), .Z(n450) );
  OR2 C9921 ( .A(n447), .B(n448), .Z(n451) );
  OR2 C9931 ( .A(n449), .B(n450), .Z(n452) );
  OR2 C997 ( .A(n5261), .B(n324), .Z(n456) );
  OR2 C998 ( .A(n325), .B(n326), .Z(n457) );
  OR2 C999 ( .A(n327), .B(n328), .Z(n458) );
  OR2 C1000 ( .A(n5270), .B(n5281), .Z(n459) );
  OR2 C10011 ( .A(n331), .B(n5284), .Z(n460) );
  OR2 C10021 ( .A(n5279), .B(n5277), .Z(n461) );
  OR2 C10031 ( .A(n335), .B(n336), .Z(n462) );
  OR2 C10041 ( .A(n456), .B(n457), .Z(n463) );
  OR2 C10051 ( .A(n458), .B(n459), .Z(n464) );
  OR2 C10061 ( .A(n460), .B(n461), .Z(n465) );
  OR2 C10071 ( .A(n462), .B(n5288), .Z(n466) );
  OR2 C1008 ( .A(n463), .B(n464), .Z(n467) );
  OR2 C1009 ( .A(n465), .B(n466), .Z(n468) );
  OR2 C10131 ( .A(n5261), .B(n324), .Z(n472) );
  OR2 C10141 ( .A(n325), .B(n326), .Z(n473) );
  OR2 C10151 ( .A(n327), .B(n328), .Z(n474) );
  OR2 C10161 ( .A(n5270), .B(n5281), .Z(n475) );
  OR2 C10171 ( .A(n331), .B(n5284), .Z(n476) );
  OR2 C10181 ( .A(n8645), .B(n334), .Z(n477) );
  OR2 C10191 ( .A(n335), .B(n336), .Z(n478) );
  OR2 C1020 ( .A(n472), .B(n473), .Z(n479) );
  OR2 C1021 ( .A(n474), .B(n475), .Z(n480) );
  OR2 C1022 ( .A(n476), .B(n477), .Z(n481) );
  OR2 C1023 ( .A(n478), .B(n5288), .Z(n482) );
  OR2 C1024 ( .A(n479), .B(n480), .Z(n483) );
  OR2 C1025 ( .A(n481), .B(n482), .Z(n484) );
  OR2 C10291 ( .A(n5261), .B(n324), .Z(n488) );
  OR2 C10301 ( .A(n325), .B(n326), .Z(n489) );
  OR2 C10311 ( .A(n327), .B(n328), .Z(n490) );
  OR2 C10321 ( .A(n5270), .B(n5281), .Z(n491) );
  OR2 C1033 ( .A(n331), .B(n8646), .Z(n492) );
  OR2 C1034 ( .A(n5279), .B(n334), .Z(n493) );
  OR2 C1035 ( .A(n335), .B(n336), .Z(n494) );
  OR2 C1036 ( .A(n488), .B(n489), .Z(n495) );
  OR2 C1037 ( .A(n490), .B(n491), .Z(n496) );
  OR2 C1038 ( .A(n492), .B(n493), .Z(n497) );
  OR2 C1039 ( .A(n494), .B(n5288), .Z(n498) );
  OR2 C1040 ( .A(n495), .B(n496), .Z(n499) );
  OR2 C10411 ( .A(n497), .B(n498), .Z(n500) );
  OR2 C10451 ( .A(n5261), .B(n324), .Z(n504) );
  OR2 C10461 ( .A(n325), .B(n326), .Z(n505) );
  OR2 C10471 ( .A(n327), .B(n328), .Z(n506) );
  OR2 C1048 ( .A(n5270), .B(n5281), .Z(n507) );
  OR2 C1049 ( .A(n5282), .B(n5284), .Z(n508) );
  OR2 C1050 ( .A(n5279), .B(n334), .Z(n509) );
  OR2 C10511 ( .A(n335), .B(n336), .Z(n510) );
  OR2 C10521 ( .A(n504), .B(n505), .Z(n511) );
  OR2 C10531 ( .A(n506), .B(n507), .Z(n512) );
  OR2 C10541 ( .A(n508), .B(n509), .Z(n513) );
  OR2 C10551 ( .A(n510), .B(n5288), .Z(n514) );
  OR2 C10561 ( .A(n511), .B(n512), .Z(n515) );
  OR2 C10571 ( .A(n513), .B(n514), .Z(n516) );
  OR2 C1061 ( .A(n5261), .B(n324), .Z(n520) );
  OR2 C1062 ( .A(n325), .B(n326), .Z(n521) );
  OR2 C1063 ( .A(n327), .B(n328), .Z(n522) );
  OR2 C1064 ( .A(n5270), .B(n8643), .Z(n523) );
  OR2 C1065 ( .A(n331), .B(n5284), .Z(n524) );
  OR2 C10661 ( .A(n5279), .B(n334), .Z(n525) );
  OR2 C10671 ( .A(n335), .B(n336), .Z(n526) );
  OR2 C10681 ( .A(n520), .B(n521), .Z(n527) );
  OR2 C10691 ( .A(n522), .B(n523), .Z(n528) );
  OR2 C10701 ( .A(n524), .B(n525), .Z(n529) );
  OR2 C10711 ( .A(n526), .B(n5288), .Z(n530) );
  OR2 C10721 ( .A(n527), .B(n528), .Z(n531) );
  OR2 C1073 ( .A(n529), .B(n530), .Z(n532) );
  OR2 C10771 ( .A(n5261), .B(n324), .Z(n536) );
  OR2 C10781 ( .A(n325), .B(n326), .Z(n537) );
  OR2 C10791 ( .A(n327), .B(n328), .Z(n538) );
  OR2 C10801 ( .A(n8642), .B(n5281), .Z(n539) );
  OR2 C10811 ( .A(n331), .B(n5284), .Z(n540) );
  OR2 C10821 ( .A(n5279), .B(n334), .Z(n541) );
  OR2 C10831 ( .A(n335), .B(n336), .Z(n542) );
  OR2 C1084 ( .A(n536), .B(n537), .Z(n543) );
  OR2 C1085 ( .A(n538), .B(n539), .Z(n544) );
  OR2 C1086 ( .A(n540), .B(n541), .Z(n545) );
  OR2 C1087 ( .A(n542), .B(n5288), .Z(n546) );
  OR2 C1088 ( .A(n543), .B(n544), .Z(n547) );
  OR2 C1089 ( .A(n545), .B(n546), .Z(n548) );
  OR2 C10931 ( .A(n5261), .B(n324), .Z(n552) );
  OR2 C10941 ( .A(n325), .B(n326), .Z(n553) );
  OR2 C10951 ( .A(n327), .B(n5269), .Z(n554) );
  OR2 C10961 ( .A(n5270), .B(n5281), .Z(n555) );
  OR2 C1097 ( .A(n331), .B(n5284), .Z(n556) );
  OR2 C1098 ( .A(n5279), .B(n334), .Z(n557) );
  OR2 C1099 ( .A(n335), .B(n336), .Z(n558) );
  OR2 C1100 ( .A(n552), .B(n553), .Z(n559) );
  OR2 C11011 ( .A(n554), .B(n555), .Z(n560) );
  OR2 C11021 ( .A(n556), .B(n557), .Z(n561) );
  OR2 C11031 ( .A(n558), .B(n5288), .Z(n562) );
  OR2 C11041 ( .A(n559), .B(n560), .Z(n563) );
  OR2 C11051 ( .A(n561), .B(n562), .Z(n564) );
  OR2 C1109 ( .A(n5261), .B(n324), .Z(n568) );
  OR2 C1110 ( .A(n325), .B(n326), .Z(n569) );
  OR2 C1111 ( .A(n5236), .B(n328), .Z(n570) );
  OR2 C1112 ( .A(n5270), .B(n5281), .Z(n571) );
  OR2 C1113 ( .A(n331), .B(n5284), .Z(n572) );
  OR2 C11141 ( .A(n5279), .B(n334), .Z(n573) );
  OR2 C11151 ( .A(n335), .B(n336), .Z(n574) );
  OR2 C11161 ( .A(n568), .B(n569), .Z(n575) );
  OR2 C11171 ( .A(n570), .B(n571), .Z(n576) );
  OR2 C11181 ( .A(n572), .B(n573), .Z(n577) );
  OR2 C11191 ( .A(n574), .B(n5288), .Z(n578) );
  OR2 C11201 ( .A(n575), .B(n576), .Z(n579) );
  OR2 C1121 ( .A(n577), .B(n578), .Z(n580) );
  OR2 C1125 ( .A(n5261), .B(n324), .Z(n584) );
  OR2 C11261 ( .A(n325), .B(n5259), .Z(n585) );
  OR2 C11271 ( .A(n327), .B(n328), .Z(n586) );
  OR2 C11281 ( .A(n5270), .B(n5281), .Z(n587) );
  OR2 C11291 ( .A(n331), .B(n5284), .Z(n588) );
  OR2 C11301 ( .A(n5279), .B(n334), .Z(n589) );
  OR2 C11311 ( .A(n335), .B(n336), .Z(n590) );
  OR2 C11321 ( .A(n584), .B(n585), .Z(n591) );
  OR2 C1133 ( .A(n586), .B(n587), .Z(n592) );
  OR2 C1134 ( .A(n588), .B(n589), .Z(n593) );
  OR2 C1135 ( .A(n590), .B(n5288), .Z(n594) );
  OR2 C1136 ( .A(n591), .B(n592), .Z(n595) );
  OR2 C1137 ( .A(n593), .B(n594), .Z(n596) );
  OR2 C11411 ( .A(n5261), .B(n324), .Z(n600) );
  OR2 C11421 ( .A(n5264), .B(n326), .Z(n601) );
  OR2 C11431 ( .A(n327), .B(n328), .Z(n602) );
  OR2 C11441 ( .A(n5270), .B(n5281), .Z(n603) );
  OR2 C11451 ( .A(n331), .B(n5284), .Z(n604) );
  OR2 C1146 ( .A(n5279), .B(n334), .Z(n605) );
  OR2 C1147 ( .A(n335), .B(n336), .Z(n606) );
  OR2 C1148 ( .A(n600), .B(n601), .Z(n607) );
  OR2 C1149 ( .A(n602), .B(n603), .Z(n608) );
  OR2 C1150 ( .A(n604), .B(n605), .Z(n609) );
  OR2 C1151 ( .A(n606), .B(n5288), .Z(n610) );
  OR2 C1152 ( .A(n607), .B(n608), .Z(n611) );
  OR2 C1153 ( .A(n609), .B(n610), .Z(n612) );
  OR2 C11571 ( .A(n5261), .B(n5263), .Z(n616) );
  OR2 C11581 ( .A(n325), .B(n326), .Z(n617) );
  OR2 C11591 ( .A(n327), .B(n328), .Z(n618) );
  OR2 C11601 ( .A(n5270), .B(n5281), .Z(n619) );
  OR2 C1161 ( .A(n331), .B(n5284), .Z(n620) );
  OR2 C1162 ( .A(n5279), .B(n334), .Z(n621) );
  OR2 C1163 ( .A(n335), .B(n336), .Z(n622) );
  OR2 C11641 ( .A(n616), .B(n617), .Z(n623) );
  OR2 C11651 ( .A(n618), .B(n619), .Z(n624) );
  OR2 C11661 ( .A(n620), .B(n621), .Z(n625) );
  OR2 C11671 ( .A(n622), .B(n5288), .Z(n626) );
  OR2 C11681 ( .A(n623), .B(n624), .Z(n627) );
  OR2 C11691 ( .A(n625), .B(n626), .Z(n628) );
  OR2 C1173 ( .A(n8641), .B(n324), .Z(n632) );
  OR2 C1174 ( .A(n325), .B(n326), .Z(n633) );
  OR2 C1175 ( .A(n327), .B(n328), .Z(n634) );
  OR2 C1176 ( .A(n5270), .B(n5281), .Z(n635) );
  OR2 C1177 ( .A(n331), .B(n5284), .Z(n636) );
  OR2 C1178 ( .A(n5279), .B(n334), .Z(n637) );
  OR2 C11791 ( .A(n335), .B(n336), .Z(n638) );
  OR2 C11801 ( .A(n632), .B(n633), .Z(n639) );
  OR2 C11811 ( .A(n634), .B(n635), .Z(n640) );
  OR2 C11821 ( .A(n636), .B(n637), .Z(n641) );
  OR2 C11831 ( .A(n638), .B(n5288), .Z(n642) );
  OR2 C11841 ( .A(n639), .B(n640), .Z(n643) );
  OR2 C11851 ( .A(n641), .B(n642), .Z(n644) );
  OR2 C19411 ( .A(n5627), .B(n5628), .Z(n1219) );
  OR2 C19421 ( .A(U4_DATA1_6), .B(n1219), .Z(n1220) );
  OR2 C19431 ( .A(U4_DATA1_5), .B(n1220), .Z(n1221) );
  OR2 C19441 ( .A(U4_DATA1_4), .B(n1221), .Z(n1222) );
  OR2 C19451 ( .A(U4_DATA1_3), .B(n1222), .Z(n1223) );
  OR2 C19461 ( .A(U4_DATA1_2), .B(n1223), .Z(n1224) );
  OR2 C19471 ( .A(U4_DATA1_1), .B(n1224), .Z(n1225) );
  OR2 C19481 ( .A(U4_DATA1_0), .B(n1225), .Z(n1226) );
  OR2 C19511 ( .A(U4_DATA1_7), .B(n5628), .Z(n1228) );
  OR2 C19521 ( .A(U4_DATA1_6), .B(n1228), .Z(n1229) );
  OR2 C19531 ( .A(U4_DATA1_5), .B(n1229), .Z(n1230) );
  OR2 C19541 ( .A(U4_DATA1_4), .B(n1230), .Z(n1231) );
  OR2 C19551 ( .A(U4_DATA1_3), .B(n1231), .Z(n1232) );
  OR2 C19561 ( .A(U4_DATA1_2), .B(n1232), .Z(n1233) );
  OR2 C19571 ( .A(U4_DATA1_1), .B(n1233), .Z(n1234) );
  OR2 C19581 ( .A(U4_DATA1_0), .B(n1234), .Z(n1235) );
  OR2 C19611 ( .A(n5627), .B(U4_DATA1_8), .Z(n1237) );
  OR2 C19621 ( .A(U4_DATA1_6), .B(n1237), .Z(n1238) );
  OR2 C19631 ( .A(U4_DATA1_5), .B(n1238), .Z(n1239) );
  OR2 C19641 ( .A(U4_DATA1_4), .B(n1239), .Z(n1240) );
  OR2 C19651 ( .A(U4_DATA1_3), .B(n1240), .Z(n1241) );
  OR2 C19661 ( .A(U4_DATA1_2), .B(n1241), .Z(n1242) );
  OR2 C19671 ( .A(U4_DATA1_1), .B(n1242), .Z(n1243) );
  OR2 C19681 ( .A(U4_DATA1_0), .B(n1243), .Z(n1244) );
  OR2 C19731 ( .A(U4_DATA1_7), .B(U4_DATA1_8), .Z(n1249) );
  OR2 C19741 ( .A(U4_DATA1_6), .B(n1249), .Z(n1250) );
  OR2 C19751 ( .A(U4_DATA1_5), .B(n1250), .Z(n1251) );
  OR2 C19761 ( .A(U4_DATA1_4), .B(n1251), .Z(n1252) );
  OR2 C19771 ( .A(U4_DATA1_3), .B(n1252), .Z(n1253) );
  OR2 C19781 ( .A(U4_DATA1_2), .B(n1253), .Z(n1254) );
  OR2 C19791 ( .A(U4_DATA1_1), .B(n1254), .Z(n1255) );
  OR2 C19801 ( .A(U4_DATA1_0), .B(n1255), .Z(n1256) );
  OR2 C19861 ( .A(n5321), .B(U157_Z_2), .Z(n1262) );
  OR2 C19871 ( .A(U156_Z_0), .B(n1262), .Z(n1263) );
  OR2 C19881 ( .A(n5319), .B(n1263), .Z(n1264) );
  OR2 C19891 ( .A(n5318), .B(n1264), .Z(n1265) );
  OR2 C19901 ( .A(n5317), .B(n1265), .Z(n1266) );
  OR2 C19911 ( .A(U158_Z_0), .B(n1266), .Z(n1267) );
  OR2 C19921 ( .A(U159_Z_0), .B(n1267), .Z(n1268) );
  OR2 C19961 ( .A(U156_Z_15), .B(U156_Z_16), .Z(n1272) );
  OR2 C19971 ( .A(U156_Z_14), .B(n1272), .Z(n1273) );
  OR2 C19981 ( .A(U156_Z_13), .B(n1273), .Z(n1274) );
  OR2 C19991 ( .A(U156_Z_12), .B(n1274), .Z(n1275) );
  OR2 C20001 ( .A(n5371), .B(n1275), .Z(n1276) );
  OR2 C20011 ( .A(n5370), .B(n1276), .Z(n1277) );
  OR2 C20021 ( .A(U158_Z_5), .B(n1277), .Z(n1278) );
  OR2 C20061 ( .A(U156_Z_10), .B(U156_Z_11), .Z(n1282) );
  OR2 C2007 ( .A(U156_Z_9), .B(n1282), .Z(n1283) );
  OR2 C20081 ( .A(U156_Z_8), .B(n1283), .Z(n1284) );
  OR2 C20091 ( .A(U156_Z_7), .B(n1284), .Z(n1285) );
  OR2 C20101 ( .A(n5353), .B(n1285), .Z(n1286) );
  OR2 C20111 ( .A(n5352), .B(n1286), .Z(n1287) );
  OR2 C20121 ( .A(U159_Z_3), .B(n1287), .Z(n1288) );
  OR2 C20161 ( .A(U156_Z_32), .B(U156_Z_33), .Z(n1292) );
  OR2 C20171 ( .A(U156_Z_31), .B(n1292), .Z(n1293) );
  OR2 C20181 ( .A(U156_Z_30), .B(n1293), .Z(n1294) );
  OR2 C20191 ( .A(U156_Z_29), .B(n1294), .Z(n1295) );
  OR2 C20201 ( .A(n5446), .B(n1295), .Z(n1296) );
  OR2 C20211 ( .A(n5445), .B(n1296), .Z(n1297) );
  OR2 C20221 ( .A(U158_Z_13), .B(n1297), .Z(n1298) );
  OR2 C2026 ( .A(U156_Z_5), .B(U156_Z_6), .Z(n1302) );
  OR2 C2027 ( .A(U156_Z_4), .B(n1302), .Z(n1303) );
  OR2 C2028 ( .A(U156_Z_3), .B(n1303), .Z(n1304) );
  OR2 C2029 ( .A(U156_Z_2), .B(n1304), .Z(n1305) );
  OR2 C2030 ( .A(n5335), .B(n1305), .Z(n1306) );
  OR2 C20311 ( .A(n5334), .B(n1306), .Z(n1307) );
  OR2 C20321 ( .A(U159_Z_2), .B(n1307), .Z(n1308) );
  OR2 C20361 ( .A(U156_Z_27), .B(U156_Z_28), .Z(n1312) );
  OR2 C2037 ( .A(U156_Z_26), .B(n1312), .Z(n1313) );
  OR2 C2038 ( .A(U156_Z_25), .B(n1313), .Z(n1314) );
  OR2 C20391 ( .A(U156_Z_24), .B(n1314), .Z(n1315) );
  OR2 C2040 ( .A(n5428), .B(n1315), .Z(n1316) );
  OR2 C20411 ( .A(n5427), .B(n1316), .Z(n1317) );
  OR2 C20421 ( .A(U159_Z_7), .B(n1317), .Z(n1318) );
  OR2 C2046 ( .A(U156_Z_1), .B(U157_Z_2), .Z(n1321) );
  OR2 C20471 ( .A(U156_Z_0), .B(n1321), .Z(n1322) );
  OR2 C20481 ( .A(U157_Z_1), .B(n1322), .Z(n1323) );
  OR2 C2049 ( .A(U157_Z_0), .B(n1323), .Z(n1324) );
  OR2 C20501 ( .A(n5317), .B(n1324), .Z(n1325) );
  OR2 C20511 ( .A(n5316), .B(n1325), .Z(n1326) );
  OR2 C20521 ( .A(U159_Z_0), .B(n1326), .Z(n1327) );
  OR2 C2056 ( .A(U156_Z_22), .B(U156_Z_23), .Z(n1331) );
  OR2 C2057 ( .A(U156_Z_21), .B(n1331), .Z(n1332) );
  OR2 C20581 ( .A(U156_Z_20), .B(n1332), .Z(n1333) );
  OR2 C20591 ( .A(U156_Z_19), .B(n1333), .Z(n1334) );
  OR2 C2060 ( .A(n5410), .B(n1334), .Z(n1335) );
  OR2 C2061 ( .A(n5409), .B(n1335), .Z(n1336) );
  OR2 C20621 ( .A(U159_Z_6), .B(n1336), .Z(n1337) );
  OR2 C2068 ( .A(n5396), .B(U157_Z_5), .Z(n1343) );
  OR2 C20691 ( .A(U156_Z_17), .B(n1343), .Z(n1344) );
  OR2 C20701 ( .A(n5394), .B(n1344), .Z(n1345) );
  OR2 C2071 ( .A(n5393), .B(n1345), .Z(n1346) );
  OR2 C2072 ( .A(n5392), .B(n1346), .Z(n1347) );
  OR2 C20731 ( .A(U158_Z_8), .B(n1347), .Z(n1348) );
  OR2 C2074 ( .A(U159_Z_4), .B(n1348), .Z(n1349) );
  OR2 C2078 ( .A(U156_Z_18), .B(U157_Z_5), .Z(n1352) );
  OR2 C2079 ( .A(U156_Z_17), .B(n1352), .Z(n1353) );
  OR2 C2080 ( .A(U157_Z_4), .B(n1353), .Z(n1354) );
  OR2 C2081 ( .A(U157_Z_3), .B(n1354), .Z(n1355) );
  OR2 C2082 ( .A(n5392), .B(n1355), .Z(n1356) );
  OR2 C2083 ( .A(n5391), .B(n1356), .Z(n1357) );
  OR2 C2084 ( .A(U159_Z_4), .B(n1357), .Z(n1358) );
  OR2 C2093 ( .A(n5375), .B(n5376), .Z(n1365) );
  OR2 C2094 ( .A(n5374), .B(n1365), .Z(n1366) );
  OR2 C2095 ( .A(n5373), .B(n1366), .Z(n1367) );
  OR2 C2096 ( .A(n5372), .B(n1367), .Z(n1368) );
  OR2 C2097 ( .A(n5371), .B(n1368), .Z(n1369) );
  OR2 C2098 ( .A(n5370), .B(n1369), .Z(n1370) );
  OR2 C2099 ( .A(U158_Z_5), .B(n1370), .Z(n1371) );
  OR2 C2108 ( .A(n5357), .B(n5358), .Z(n1378) );
  OR2 C2109 ( .A(n5356), .B(n1378), .Z(n1379) );
  OR2 C2110 ( .A(n5355), .B(n1379), .Z(n1380) );
  OR2 C21111 ( .A(n5354), .B(n1380), .Z(n1381) );
  OR2 C2112 ( .A(n5353), .B(n1381), .Z(n1382) );
  OR2 C2113 ( .A(n5352), .B(n1382), .Z(n1383) );
  OR2 C2114 ( .A(U159_Z_3), .B(n1383), .Z(n1384) );
  OR2 C2123 ( .A(n5450), .B(n5451), .Z(n1391) );
  OR2 C2124 ( .A(n5449), .B(n1391), .Z(n1392) );
  OR2 C2125 ( .A(n5448), .B(n1392), .Z(n1393) );
  OR2 C2126 ( .A(n5447), .B(n1393), .Z(n1394) );
  OR2 C2127 ( .A(n5446), .B(n1394), .Z(n1395) );
  OR2 C2128 ( .A(n5445), .B(n1395), .Z(n1396) );
  OR2 C2129 ( .A(U158_Z_13), .B(n1396), .Z(n1397) );
  OR2 C2138 ( .A(n5339), .B(n5340), .Z(n1404) );
  OR2 C2139 ( .A(n5338), .B(n1404), .Z(n1405) );
  OR2 C2140 ( .A(n5337), .B(n1405), .Z(n1406) );
  OR2 C2141 ( .A(n5336), .B(n1406), .Z(n1407) );
  OR2 C2142 ( .A(n5335), .B(n1407), .Z(n1408) );
  OR2 C2143 ( .A(n5334), .B(n1408), .Z(n1409) );
  OR2 C2144 ( .A(U159_Z_2), .B(n1409), .Z(n1410) );
  OR2 C2153 ( .A(n5432), .B(n5433), .Z(n1417) );
  OR2 C2154 ( .A(n5431), .B(n1417), .Z(n1418) );
  OR2 C2155 ( .A(n5430), .B(n1418), .Z(n1419) );
  OR2 C2156 ( .A(n5429), .B(n1419), .Z(n1420) );
  OR2 C2157 ( .A(n5428), .B(n1420), .Z(n1421) );
  OR2 C2158 ( .A(n5427), .B(n1421), .Z(n1422) );
  OR2 C2159 ( .A(U159_Z_7), .B(n1422), .Z(n1423) );
  OR2 C2168 ( .A(n5321), .B(n5322), .Z(n1427) );
  OR2 C2169 ( .A(n5320), .B(n1427), .Z(n1428) );
  OR2 C2170 ( .A(n5319), .B(n1428), .Z(n1429) );
  OR2 C21711 ( .A(n5318), .B(n1429), .Z(n1430) );
  OR2 C2172 ( .A(n5317), .B(n1430), .Z(n1431) );
  OR2 C2173 ( .A(n5316), .B(n1431), .Z(n1432) );
  OR2 C2174 ( .A(U159_Z_0), .B(n1432), .Z(n1433) );
  OR2 C2183 ( .A(n5414), .B(n5415), .Z(n1440) );
  OR2 C2184 ( .A(n5413), .B(n1440), .Z(n1441) );
  OR2 C2185 ( .A(n5412), .B(n1441), .Z(n1442) );
  OR2 C2186 ( .A(n5411), .B(n1442), .Z(n1443) );
  OR2 C2187 ( .A(n5410), .B(n1443), .Z(n1444) );
  OR2 C2188 ( .A(n5409), .B(n1444), .Z(n1445) );
  OR2 C2189 ( .A(U159_Z_6), .B(n1445), .Z(n1446) );
  OR2 C2198 ( .A(n5396), .B(n5397), .Z(n1450) );
  OR2 C2199 ( .A(n5395), .B(n1450), .Z(n1451) );
  OR2 C2200 ( .A(n5394), .B(n1451), .Z(n1452) );
  OR2 C2201 ( .A(n5393), .B(n1452), .Z(n1453) );
  OR2 C2202 ( .A(n5392), .B(n1453), .Z(n1454) );
  OR2 C2203 ( .A(n5391), .B(n1454), .Z(n1455) );
  OR2 C2204 ( .A(U159_Z_4), .B(n1455), .Z(n1456) );
  OR2 C2216 ( .A(U156_Z_12), .B(n1367), .Z(n1459) );
  OR2 C2217 ( .A(n5371), .B(n1459), .Z(n1460) );
  OR2 C2218 ( .A(n5370), .B(n1460), .Z(n1461) );
  OR2 C2219 ( .A(n5362), .B(n1461), .Z(n1462) );
  OR2 C2231 ( .A(U156_Z_7), .B(n1380), .Z(n1465) );
  OR2 C2232 ( .A(n5353), .B(n1465), .Z(n1466) );
  OR2 C2233 ( .A(n5352), .B(n1466), .Z(n1467) );
  OR2 C2234 ( .A(n5344), .B(n1467), .Z(n1468) );
  OR2 C2246 ( .A(U156_Z_29), .B(n1393), .Z(n1471) );
  OR2 C2247 ( .A(n5446), .B(n1471), .Z(n1472) );
  OR2 C2248 ( .A(n5445), .B(n1472), .Z(n1473) );
  OR2 C2249 ( .A(n5437), .B(n1473), .Z(n1474) );
  OR2 C2261 ( .A(U156_Z_2), .B(n1406), .Z(n1477) );
  OR2 C2262 ( .A(n5335), .B(n1477), .Z(n1478) );
  OR2 C2263 ( .A(n5334), .B(n1478), .Z(n1479) );
  OR2 C2264 ( .A(n5326), .B(n1479), .Z(n1480) );
  OR2 C2276 ( .A(U156_Z_24), .B(n1419), .Z(n1483) );
  OR2 C2277 ( .A(n5428), .B(n1483), .Z(n1484) );
  OR2 C2278 ( .A(n5427), .B(n1484), .Z(n1485) );
  OR2 C2279 ( .A(n5419), .B(n1485), .Z(n1486) );
  OR2 C2291 ( .A(U157_Z_0), .B(n1429), .Z(n1489) );
  OR2 C2292 ( .A(n5317), .B(n1489), .Z(n1490) );
  OR2 C2293 ( .A(n5316), .B(n1490), .Z(n1491) );
  OR2 C2294 ( .A(n5306), .B(n1491), .Z(n1492) );
  OR2 C2306 ( .A(U156_Z_19), .B(n1442), .Z(n1495) );
  OR2 C2307 ( .A(n5410), .B(n1495), .Z(n1496) );
  OR2 C2308 ( .A(n5409), .B(n1496), .Z(n1497) );
  OR2 C2309 ( .A(n5401), .B(n1497), .Z(n1498) );
  OR2 C2311 ( .A(U154_Z_4), .B(U154_Z_5), .Z(n1500) );
  OR2 C2312 ( .A(U154_Z_3), .B(n1500), .Z(n1501) );
  OR2 C2313 ( .A(U155_Z_1), .B(n1501), .Z(n1502) );
  OR2 C2314 ( .A(U154_Z_2), .B(n1502), .Z(n1503) );
  OR2 C2315 ( .A(U154_Z_1), .B(n1503), .Z(n1504) );
  OR2 C2316 ( .A(U154_Z_0), .B(n1504), .Z(n1505) );
  OR2 C2317 ( .A(U155_Z_0), .B(n1505), .Z(n1506) );
  OR2 C2329 ( .A(U157_Z_3), .B(n1452), .Z(n1509) );
  OR2 C2330 ( .A(n5392), .B(n1509), .Z(n1510) );
  OR2 C2331 ( .A(n5391), .B(n1510), .Z(n1511) );
  OR2 C2332 ( .A(n5381), .B(n1511), .Z(n1512) );
  OR2 C2340 ( .A(U156_Z_14), .B(n1365), .Z(n1514) );
  OR2 C2341 ( .A(n5373), .B(n1514), .Z(n1515) );
  OR2 C2342 ( .A(n5372), .B(n1515), .Z(n1516) );
  OR2 C2343 ( .A(n5371), .B(n1516), .Z(n1517) );
  OR2 C2344 ( .A(U158_Z_6), .B(n1517), .Z(n1518) );
  OR2 C2345 ( .A(U158_Z_5), .B(n1518), .Z(n1519) );
  OR2 C2353 ( .A(U156_Z_9), .B(n1378), .Z(n1521) );
  OR2 C2354 ( .A(n5355), .B(n1521), .Z(n1522) );
  OR2 C2355 ( .A(n5354), .B(n1522), .Z(n1523) );
  OR2 C2356 ( .A(n5353), .B(n1523), .Z(n1524) );
  OR2 C2357 ( .A(U158_Z_3), .B(n1524), .Z(n1525) );
  OR2 C2358 ( .A(U159_Z_3), .B(n1525), .Z(n1526) );
  OR2 C2366 ( .A(U156_Z_31), .B(n1391), .Z(n1528) );
  OR2 C2367 ( .A(n5448), .B(n1528), .Z(n1529) );
  OR2 C2368 ( .A(n5447), .B(n1529), .Z(n1530) );
  OR2 C2369 ( .A(n5446), .B(n1530), .Z(n1531) );
  OR2 C2370 ( .A(U158_Z_14), .B(n1531), .Z(n1532) );
  OR2 C2371 ( .A(U158_Z_13), .B(n1532), .Z(n1533) );
  OR2 C2379 ( .A(U156_Z_4), .B(n1404), .Z(n1535) );
  OR2 C2380 ( .A(n5337), .B(n1535), .Z(n1536) );
  OR2 C2381 ( .A(n5336), .B(n1536), .Z(n1537) );
  OR2 C2382 ( .A(n5335), .B(n1537), .Z(n1538) );
  OR2 C2383 ( .A(U158_Z_1), .B(n1538), .Z(n1539) );
  OR2 C2384 ( .A(U159_Z_2), .B(n1539), .Z(n1540) );
  OR2 C2392 ( .A(U156_Z_26), .B(n1417), .Z(n1542) );
  OR2 C2393 ( .A(n5430), .B(n1542), .Z(n1543) );
  OR2 C2394 ( .A(n5429), .B(n1543), .Z(n1544) );
  OR2 C2395 ( .A(n5428), .B(n1544), .Z(n1545) );
  OR2 C2396 ( .A(U158_Z_11), .B(n1545), .Z(n1546) );
  OR2 C2397 ( .A(U159_Z_7), .B(n1546), .Z(n1547) );
  OR2 C2405 ( .A(U156_Z_0), .B(n1427), .Z(n1549) );
  OR2 C2406 ( .A(n5319), .B(n1549), .Z(n1550) );
  OR2 C2407 ( .A(n5318), .B(n1550), .Z(n1551) );
  OR2 C2408 ( .A(n5317), .B(n1551), .Z(n1552) );
  OR2 C2409 ( .A(U158_Z_0), .B(n1552), .Z(n1553) );
  OR2 C2410 ( .A(U159_Z_0), .B(n1553), .Z(n1554) );
  OR2 C2418 ( .A(U156_Z_21), .B(n1440), .Z(n1556) );
  OR2 C2419 ( .A(n5412), .B(n1556), .Z(n1557) );
  OR2 C2420 ( .A(n5411), .B(n1557), .Z(n1558) );
  OR2 C2421 ( .A(n5410), .B(n1558), .Z(n1559) );
  OR2 C2422 ( .A(U158_Z_9), .B(n1559), .Z(n1560) );
  OR2 C2423 ( .A(U159_Z_6), .B(n1560), .Z(n1561) );
  OR2 C2431 ( .A(U156_Z_17), .B(n1450), .Z(n1563) );
  OR2 C2432 ( .A(n5394), .B(n1563), .Z(n1564) );
  OR2 C2433 ( .A(n5393), .B(n1564), .Z(n1565) );
  OR2 C2434 ( .A(n5392), .B(n1565), .Z(n1566) );
  OR2 C2435 ( .A(U158_Z_8), .B(n1566), .Z(n1567) );
  OR2 C2436 ( .A(U159_Z_4), .B(n1567), .Z(n1568) );
  OR2 C2443 ( .A(n5374), .B(n1272), .Z(n1570) );
  OR2 C2444 ( .A(n5373), .B(n1570), .Z(n1571) );
  OR2 C2445 ( .A(n5372), .B(n1571), .Z(n1572) );
  OR2 C2446 ( .A(n5371), .B(n1572), .Z(n1573) );
  OR2 C2447 ( .A(U158_Z_6), .B(n1573), .Z(n1574) );
  OR2 C2448 ( .A(U158_Z_5), .B(n1574), .Z(n1575) );
  OR2 C2455 ( .A(n5356), .B(n1282), .Z(n1577) );
  OR2 C2456 ( .A(n5355), .B(n1577), .Z(n1578) );
  OR2 C2457 ( .A(n5354), .B(n1578), .Z(n1579) );
  OR2 C2458 ( .A(n5353), .B(n1579), .Z(n1580) );
  OR2 C2459 ( .A(U158_Z_3), .B(n1580), .Z(n1581) );
  OR2 C2460 ( .A(U159_Z_3), .B(n1581), .Z(n1582) );
  OR2 C2467 ( .A(n5449), .B(n1292), .Z(n1584) );
  OR2 C2468 ( .A(n5448), .B(n1584), .Z(n1585) );
  OR2 C2469 ( .A(n5447), .B(n1585), .Z(n1586) );
  OR2 C2470 ( .A(n5446), .B(n1586), .Z(n1587) );
  OR2 C2471 ( .A(U158_Z_14), .B(n1587), .Z(n1588) );
  OR2 C2472 ( .A(U158_Z_13), .B(n1588), .Z(n1589) );
  OR2 C2479 ( .A(n5338), .B(n1302), .Z(n1591) );
  OR2 C2480 ( .A(n5337), .B(n1591), .Z(n1592) );
  OR2 C2481 ( .A(n5336), .B(n1592), .Z(n1593) );
  OR2 C2482 ( .A(n5335), .B(n1593), .Z(n1594) );
  OR2 C2483 ( .A(U158_Z_1), .B(n1594), .Z(n1595) );
  OR2 C2484 ( .A(U159_Z_2), .B(n1595), .Z(n1596) );
  OR2 C2491 ( .A(n5431), .B(n1312), .Z(n1598) );
  OR2 C2492 ( .A(n5430), .B(n1598), .Z(n1599) );
  OR2 C2493 ( .A(n5429), .B(n1599), .Z(n1600) );
  OR2 C2494 ( .A(n5428), .B(n1600), .Z(n1601) );
  OR2 C2495 ( .A(U158_Z_11), .B(n1601), .Z(n1602) );
  OR2 C2496 ( .A(U159_Z_7), .B(n1602), .Z(n1603) );
  OR2 C2503 ( .A(n5320), .B(n1321), .Z(n1605) );
  OR2 C2504 ( .A(n5319), .B(n1605), .Z(n1606) );
  OR2 C2505 ( .A(n5318), .B(n1606), .Z(n1607) );
  OR2 C2506 ( .A(n5317), .B(n1607), .Z(n1608) );
  OR2 C2507 ( .A(U158_Z_0), .B(n1608), .Z(n1609) );
  OR2 C2508 ( .A(U159_Z_0), .B(n1609), .Z(n1610) );
  OR2 C2515 ( .A(n5413), .B(n1331), .Z(n1612) );
  OR2 C2516 ( .A(n5412), .B(n1612), .Z(n1613) );
  OR2 C2517 ( .A(n5411), .B(n1613), .Z(n1614) );
  OR2 C2518 ( .A(n5410), .B(n1614), .Z(n1615) );
  OR2 C2519 ( .A(U158_Z_9), .B(n1615), .Z(n1616) );
  OR2 C2520 ( .A(U159_Z_6), .B(n1616), .Z(n1617) );
  OR2 C2527 ( .A(n5395), .B(n1352), .Z(n1619) );
  OR2 C2528 ( .A(n5394), .B(n1619), .Z(n1620) );
  OR2 C2529 ( .A(n5393), .B(n1620), .Z(n1621) );
  OR2 C2530 ( .A(n5392), .B(n1621), .Z(n1622) );
  OR2 C2531 ( .A(U158_Z_8), .B(n1622), .Z(n1623) );
  OR2 C2532 ( .A(U159_Z_4), .B(n1623), .Z(n1624) );
  OR2 C2539 ( .A(n5373), .B(n1273), .Z(n1626) );
  OR2 C2540 ( .A(n5372), .B(n1626), .Z(n1627) );
  OR2 C2541 ( .A(n5371), .B(n1627), .Z(n1628) );
  OR2 C2542 ( .A(U158_Z_6), .B(n1628), .Z(n1629) );
  OR2 C2543 ( .A(U158_Z_5), .B(n1629), .Z(n1630) );
  OR2 C2550 ( .A(n5355), .B(n1283), .Z(n1632) );
  OR2 C2551 ( .A(n5354), .B(n1632), .Z(n1633) );
  OR2 C2552 ( .A(n5353), .B(n1633), .Z(n1634) );
  OR2 C2553 ( .A(U158_Z_3), .B(n1634), .Z(n1635) );
  OR2 C2554 ( .A(U159_Z_3), .B(n1635), .Z(n1636) );
  OR2 C2561 ( .A(n5448), .B(n1293), .Z(n1638) );
  OR2 C2562 ( .A(n5447), .B(n1638), .Z(n1639) );
  OR2 C2563 ( .A(n5446), .B(n1639), .Z(n1640) );
  OR2 C2564 ( .A(U158_Z_14), .B(n1640), .Z(n1641) );
  OR2 C2565 ( .A(U158_Z_13), .B(n1641), .Z(n1642) );
  OR2 C2572 ( .A(n5337), .B(n1303), .Z(n1644) );
  OR2 C2573 ( .A(n5336), .B(n1644), .Z(n1645) );
  OR2 C2574 ( .A(n5335), .B(n1645), .Z(n1646) );
  OR2 C2575 ( .A(U158_Z_1), .B(n1646), .Z(n1647) );
  OR2 C2576 ( .A(U159_Z_2), .B(n1647), .Z(n1648) );
  OR2 C2583 ( .A(n5430), .B(n1313), .Z(n1650) );
  OR2 C2584 ( .A(n5429), .B(n1650), .Z(n1651) );
  OR2 C2585 ( .A(n5428), .B(n1651), .Z(n1652) );
  OR2 C2586 ( .A(U158_Z_11), .B(n1652), .Z(n1653) );
  OR2 C2587 ( .A(U159_Z_7), .B(n1653), .Z(n1654) );
  OR2 C2594 ( .A(n5319), .B(n1322), .Z(n1656) );
  OR2 C2595 ( .A(n5318), .B(n1656), .Z(n1657) );
  OR2 C2596 ( .A(n5317), .B(n1657), .Z(n1658) );
  OR2 C2597 ( .A(U158_Z_0), .B(n1658), .Z(n1659) );
  OR2 C2598 ( .A(U159_Z_0), .B(n1659), .Z(n1660) );
  OR2 C2605 ( .A(n5412), .B(n1332), .Z(n1662) );
  OR2 C2606 ( .A(n5411), .B(n1662), .Z(n1663) );
  OR2 C2607 ( .A(n5410), .B(n1663), .Z(n1664) );
  OR2 C2608 ( .A(U158_Z_9), .B(n1664), .Z(n1665) );
  OR2 C2609 ( .A(U159_Z_6), .B(n1665), .Z(n1666) );
  OR2 C2616 ( .A(n5394), .B(n1353), .Z(n1668) );
  OR2 C2617 ( .A(n5393), .B(n1668), .Z(n1669) );
  OR2 C2618 ( .A(n5392), .B(n1669), .Z(n1670) );
  OR2 C2619 ( .A(U158_Z_8), .B(n1670), .Z(n1671) );
  OR2 C2620 ( .A(U159_Z_4), .B(n1671), .Z(n1672) );
  OR2 C2627 ( .A(U156_Z_15), .B(n5376), .Z(n1674) );
  OR2 C2628 ( .A(n5374), .B(n1674), .Z(n1675) );
  OR2 C2629 ( .A(n5373), .B(n1675), .Z(n1676) );
  OR2 C2630 ( .A(n5372), .B(n1676), .Z(n1677) );
  OR2 C2631 ( .A(n5371), .B(n1677), .Z(n1678) );
  OR2 C2632 ( .A(U158_Z_6), .B(n1678), .Z(n1679) );
  OR2 C2633 ( .A(U158_Z_5), .B(n1679), .Z(n1680) );
  OR2 C2640 ( .A(U156_Z_10), .B(n5358), .Z(n1682) );
  OR2 C2641 ( .A(n5356), .B(n1682), .Z(n1683) );
  OR2 C2642 ( .A(n5355), .B(n1683), .Z(n1684) );
  OR2 C2643 ( .A(n5354), .B(n1684), .Z(n1685) );
  OR2 C2644 ( .A(n5353), .B(n1685), .Z(n1686) );
  OR2 C2645 ( .A(U158_Z_3), .B(n1686), .Z(n1687) );
  OR2 C2646 ( .A(U159_Z_3), .B(n1687), .Z(n1688) );
  OR2 C2653 ( .A(U156_Z_32), .B(n5451), .Z(n1690) );
  OR2 C2654 ( .A(n5449), .B(n1690), .Z(n1691) );
  OR2 C2655 ( .A(n5448), .B(n1691), .Z(n1692) );
  OR2 C2656 ( .A(n5447), .B(n1692), .Z(n1693) );
  OR2 C2657 ( .A(n5446), .B(n1693), .Z(n1694) );
  OR2 C2658 ( .A(U158_Z_14), .B(n1694), .Z(n1695) );
  OR2 C2659 ( .A(U158_Z_13), .B(n1695), .Z(n1696) );
  OR2 C2666 ( .A(U156_Z_5), .B(n5340), .Z(n1698) );
  OR2 C2667 ( .A(n5338), .B(n1698), .Z(n1699) );
  OR2 C2668 ( .A(n5337), .B(n1699), .Z(n1700) );
  OR2 C2669 ( .A(n5336), .B(n1700), .Z(n1701) );
  OR2 C2670 ( .A(n5335), .B(n1701), .Z(n1702) );
  OR2 C2671 ( .A(U158_Z_1), .B(n1702), .Z(n1703) );
  OR2 C2672 ( .A(U159_Z_2), .B(n1703), .Z(n1704) );
  OR2 C2679 ( .A(U156_Z_27), .B(n5433), .Z(n1706) );
  OR2 C2680 ( .A(n5431), .B(n1706), .Z(n1707) );
  OR2 C2681 ( .A(n5430), .B(n1707), .Z(n1708) );
  OR2 C2682 ( .A(n5429), .B(n1708), .Z(n1709) );
  OR2 C2683 ( .A(n5428), .B(n1709), .Z(n1710) );
  OR2 C2684 ( .A(U158_Z_11), .B(n1710), .Z(n1711) );
  OR2 C2685 ( .A(U159_Z_7), .B(n1711), .Z(n1712) );
  OR2 C2692 ( .A(U156_Z_1), .B(n5322), .Z(n1714) );
  OR2 C2693 ( .A(n5320), .B(n1714), .Z(n1715) );
  OR2 C2694 ( .A(n5319), .B(n1715), .Z(n1716) );
  OR2 C2695 ( .A(n5318), .B(n1716), .Z(n1717) );
  OR2 C2696 ( .A(n5317), .B(n1717), .Z(n1718) );
  OR2 C2697 ( .A(U158_Z_0), .B(n1718), .Z(n1719) );
  OR2 C2698 ( .A(U159_Z_0), .B(n1719), .Z(n1720) );
  OR2 C2705 ( .A(U156_Z_22), .B(n5415), .Z(n1722) );
  OR2 C2706 ( .A(n5413), .B(n1722), .Z(n1723) );
  OR2 C2707 ( .A(n5412), .B(n1723), .Z(n1724) );
  OR2 C2708 ( .A(n5411), .B(n1724), .Z(n1725) );
  OR2 C2709 ( .A(n5410), .B(n1725), .Z(n1726) );
  OR2 C2710 ( .A(U158_Z_9), .B(n1726), .Z(n1727) );
  OR2 C27111 ( .A(U159_Z_6), .B(n1727), .Z(n1728) );
  OR2 C2718 ( .A(U156_Z_18), .B(n5397), .Z(n1730) );
  OR2 C2719 ( .A(n5395), .B(n1730), .Z(n1731) );
  OR2 C2720 ( .A(n5394), .B(n1731), .Z(n1732) );
  OR2 C2721 ( .A(n5393), .B(n1732), .Z(n1733) );
  OR2 C2722 ( .A(n5392), .B(n1733), .Z(n1734) );
  OR2 C2723 ( .A(U158_Z_8), .B(n1734), .Z(n1735) );
  OR2 C2724 ( .A(U159_Z_4), .B(n1735), .Z(n1736) );
  OR2 C2731 ( .A(n5375), .B(U156_Z_16), .Z(n1738) );
  OR2 C2732 ( .A(n5374), .B(n1738), .Z(n1739) );
  OR2 C2733 ( .A(n5373), .B(n1739), .Z(n1740) );
  OR2 C2734 ( .A(n5372), .B(n1740), .Z(n1741) );
  OR2 C2735 ( .A(n5371), .B(n1741), .Z(n1742) );
  OR2 C2736 ( .A(U158_Z_6), .B(n1742), .Z(n1743) );
  OR2 C2737 ( .A(U158_Z_5), .B(n1743), .Z(n1744) );
  OR2 C2744 ( .A(n5357), .B(U156_Z_11), .Z(n1746) );
  OR2 C2745 ( .A(n5356), .B(n1746), .Z(n1747) );
  OR2 C2746 ( .A(n5355), .B(n1747), .Z(n1748) );
  OR2 C2747 ( .A(n5354), .B(n1748), .Z(n1749) );
  OR2 C2748 ( .A(n5353), .B(n1749), .Z(n1750) );
  OR2 C2749 ( .A(U158_Z_3), .B(n1750), .Z(n1751) );
  OR2 C2750 ( .A(U159_Z_3), .B(n1751), .Z(n1752) );
  OR2 C2757 ( .A(n5450), .B(U156_Z_33), .Z(n1754) );
  OR2 C2758 ( .A(n5449), .B(n1754), .Z(n1755) );
  OR2 C2759 ( .A(n5448), .B(n1755), .Z(n1756) );
  OR2 C2760 ( .A(n5447), .B(n1756), .Z(n1757) );
  OR2 C2761 ( .A(n5446), .B(n1757), .Z(n1758) );
  OR2 C2762 ( .A(U158_Z_14), .B(n1758), .Z(n1759) );
  OR2 C2763 ( .A(U158_Z_13), .B(n1759), .Z(n1760) );
  OR2 C2770 ( .A(n5339), .B(U156_Z_6), .Z(n1762) );
  OR2 C2771 ( .A(n5338), .B(n1762), .Z(n1763) );
  OR2 C2772 ( .A(n5337), .B(n1763), .Z(n1764) );
  OR2 C2773 ( .A(n5336), .B(n1764), .Z(n1765) );
  OR2 C2774 ( .A(n5335), .B(n1765), .Z(n1766) );
  OR2 C2775 ( .A(U158_Z_1), .B(n1766), .Z(n1767) );
  OR2 C2776 ( .A(U159_Z_2), .B(n1767), .Z(n1768) );
  OR2 C2783 ( .A(n5432), .B(U156_Z_28), .Z(n1770) );
  OR2 C2784 ( .A(n5431), .B(n1770), .Z(n1771) );
  OR2 C2785 ( .A(n5430), .B(n1771), .Z(n1772) );
  OR2 C2786 ( .A(n5429), .B(n1772), .Z(n1773) );
  OR2 C2787 ( .A(n5428), .B(n1773), .Z(n1774) );
  OR2 C2788 ( .A(U158_Z_11), .B(n1774), .Z(n1775) );
  OR2 C2789 ( .A(U159_Z_7), .B(n1775), .Z(n1776) );
  OR2 C2797 ( .A(n5320), .B(n1262), .Z(n1778) );
  OR2 C2798 ( .A(n5319), .B(n1778), .Z(n1779) );
  OR2 C2799 ( .A(n5318), .B(n1779), .Z(n1780) );
  OR2 C2800 ( .A(n5317), .B(n1780), .Z(n1781) );
  OR2 C2801 ( .A(U158_Z_0), .B(n1781), .Z(n1782) );
  OR2 C2802 ( .A(U159_Z_0), .B(n1782), .Z(n1783) );
  OR2 C2809 ( .A(n5414), .B(U156_Z_23), .Z(n1785) );
  OR2 C2810 ( .A(n5413), .B(n1785), .Z(n1786) );
  OR2 C2811 ( .A(n5412), .B(n1786), .Z(n1787) );
  OR2 C2812 ( .A(n5411), .B(n1787), .Z(n1788) );
  OR2 C2813 ( .A(n5410), .B(n1788), .Z(n1789) );
  OR2 C2814 ( .A(U158_Z_9), .B(n1789), .Z(n1790) );
  OR2 C2815 ( .A(U159_Z_6), .B(n1790), .Z(n1791) );
  OR2 C2823 ( .A(n5395), .B(n1343), .Z(n1793) );
  OR2 C2824 ( .A(n5394), .B(n1793), .Z(n1794) );
  OR2 C2825 ( .A(n5393), .B(n1794), .Z(n1795) );
  OR2 C2826 ( .A(n5392), .B(n1795), .Z(n1796) );
  OR2 C2827 ( .A(U158_Z_8), .B(n1796), .Z(n1797) );
  OR2 C2828 ( .A(U159_Z_4), .B(n1797), .Z(n1798) );
  OR2 C2839 ( .A(n5362), .B(n1277), .Z(n1800) );
  OR2 C2851 ( .A(n5344), .B(n1287), .Z(n1803) );
  OR2 C2863 ( .A(n5437), .B(n1297), .Z(n1806) );
  OR2 C2875 ( .A(n5326), .B(n1307), .Z(n1809) );
  OR2 C2887 ( .A(n5419), .B(n1317), .Z(n1812) );
  OR2 C2899 ( .A(n5306), .B(n1326), .Z(n1815) );
  OR2 C2911 ( .A(n5401), .B(n1336), .Z(n1818) );
  OR2 C2923 ( .A(n5381), .B(n1357), .Z(n1821) );
  OR2 C2938 ( .A(U158_Z_14), .B(n1395), .Z(n1824) );
  OR2 C2939 ( .A(n5437), .B(n1824), .Z(n1825) );
  OR2 C2953 ( .A(U158_Z_11), .B(n1421), .Z(n1827) );
  OR2 C2954 ( .A(n5419), .B(n1827), .Z(n1828) );
  OR2 C2968 ( .A(U158_Z_9), .B(n1444), .Z(n1830) );
  OR2 C2969 ( .A(n5401), .B(n1830), .Z(n1831) );
  OR2 C2983 ( .A(U158_Z_8), .B(n1454), .Z(n1833) );
  OR2 C2984 ( .A(n5381), .B(n1833), .Z(n1834) );
  OR2 C2998 ( .A(U158_Z_6), .B(n1369), .Z(n1836) );
  OR2 C2999 ( .A(n5362), .B(n1836), .Z(n1837) );
  OR2 C3013 ( .A(U158_Z_3), .B(n1382), .Z(n1839) );
  OR2 C3014 ( .A(n5344), .B(n1839), .Z(n1840) );
  OR2 C3028 ( .A(U158_Z_1), .B(n1408), .Z(n1842) );
  OR2 C3029 ( .A(n5326), .B(n1842), .Z(n1843) );
  OR2 C3043 ( .A(U158_Z_0), .B(n1431), .Z(n1845) );
  OR2 C3044 ( .A(n5306), .B(n1845), .Z(n1846) );
  OR2 C3057 ( .A(U159_Z_1), .B(n1430), .Z(n1848) );
  OR2 C3058 ( .A(n5316), .B(n1848), .Z(n1849) );
  OR2 C3059 ( .A(n5306), .B(n1849), .Z(n1850) );
  OR2 C3066 ( .A(U156_Z_0), .B(n1714), .Z(n1852) );
  OR2 C3067 ( .A(n5319), .B(n1852), .Z(n1853) );
  OR2 C3068 ( .A(n5318), .B(n1853), .Z(n1854) );
  OR2 C3069 ( .A(n5317), .B(n1854), .Z(n1855) );
  OR2 C3070 ( .A(U158_Z_0), .B(n1855), .Z(n1856) );
  OR2 C3071 ( .A(U159_Z_0), .B(n1856), .Z(n1857) );
  OR2 C3096 ( .A(U159_Z_5), .B(n1453), .Z(n1859) );
  OR2 C3097 ( .A(n5391), .B(n1859), .Z(n1860) );
  OR2 C3098 ( .A(n5381), .B(n1860), .Z(n1861) );
  OR2 C3105 ( .A(U156_Z_17), .B(n1730), .Z(n1863) );
  OR2 C3106 ( .A(n5394), .B(n1863), .Z(n1864) );
  OR2 C3107 ( .A(n5393), .B(n1864), .Z(n1865) );
  OR2 C3108 ( .A(n5392), .B(n1865), .Z(n1866) );
  OR2 C3109 ( .A(U158_Z_8), .B(n1866), .Z(n1867) );
  OR2 C3110 ( .A(U159_Z_4), .B(n1867), .Z(n1868) );
  OR2 C5223 ( .A(n1870), .B(n127), .Z(U59_DATA1_0) );
  OR2 C5227 ( .A(n1871), .B(n127), .Z(U59_DATA1_1) );
  OR2 C5254 ( .A(n1872), .B(n143), .Z(U57_DATA1_0) );
  OR2 C5258 ( .A(n1873), .B(n143), .Z(U57_DATA1_1) );
  OR2 C5285 ( .A(n1874), .B(n159), .Z(U55_DATA1_1) );
  OR2 C5289 ( .A(n1875), .B(n159), .Z(U54_DATA1_0) );
  OR2 C5316 ( .A(n1876), .B(n175), .Z(U52_DATA1_1) );
  OR2 C5320 ( .A(n1877), .B(n175), .Z(U52_DATA1_2) );
  OR2 C5347 ( .A(n1878), .B(n191), .Z(U61_DATA2_1) );
  OR2 C53511 ( .A(n1879), .B(n191), .Z(U61_DATA2_2) );
  OR2 C5378 ( .A(n1880), .B(n207), .Z(U61_DATA2_8) );
  OR2 C5382 ( .A(n1881), .B(n207), .Z(U61_DATA2_9) );
  OR2 C5409 ( .A(n1882), .B(n223), .Z(U61_DATA2_15) );
  OR2 C5413 ( .A(n1883), .B(n223), .Z(U61_DATA2_16) );
  OR2 C5440 ( .A(n1884), .B(n239), .Z(U61_DATA2_22) );
  OR2 C5444 ( .A(n1885), .B(n239), .Z(U61_DATA2_23) );
  OR2 C5528 ( .A(n338), .B(n339), .Z(n327) );
  OR2 C5559 ( .A(n1886), .B(n1887), .Z(U40_DATA2_0) );
  OR2 C5563 ( .A(n1888), .B(n1889), .Z(U40_DATA2_1) );
  OR2 C5570 ( .A(n1890), .B(n1891), .Z(U40_DATA2_2) );
  OR2 C5577 ( .A(n1892), .B(n1893), .Z(U40_DATA2_3) );
  OR2 C5584 ( .A(n1894), .B(n1895), .Z(U40_DATA2_4) );
  OR2 C5594 ( .A(n1896), .B(n1897), .Z(U40_DATA2_5) );
  OR2 C5601 ( .A(n1899), .B(n1900), .Z(U40_DATA2_6) );
  OR2 C5608 ( .A(n1901), .B(n1900), .Z(U40_DATA2_7) );
  OR2 C5614 ( .A(n5246), .B(n5245), .Z(n1906) );
  OR2 C5615 ( .A(n1905), .B(n1906), .Z(n1907) );
  OR2 C5664 ( .A(n1909), .B(n5245), .Z(n1910) );
  OR2 C5726 ( .A(n1898), .B(n5249), .Z(n1914) );
  OR2 C5763 ( .A(n5257), .B(n5254), .Z(n1919) );
  OR2 C5797 ( .A(n1918), .B(n5248), .Z(n1924) );
  OR2 C5834 ( .A(n5248), .B(n5247), .Z(n1926) );
  OR2 C5835 ( .A(n1918), .B(n1926), .Z(n1927) );
  OR2 C5877 ( .A(n1918), .B(n1929), .Z(n1930) );
  OR2 C5911 ( .A(n816), .B(n817), .Z(n1932) );
  OR2 C5914 ( .A(n816), .B(n750), .Z(n1934) );
  OR2 C6102 ( .A(n1115), .B(n940), .Z(n1935) );
  AN2 C6252 ( .A(n5684), .B(n5294), .Z(n99) );
  AN2 C6263 ( .A(n1947), .B(n1327), .Z(n110) );
  AN2 C6264 ( .A(n1946), .B(n1433), .Z(n1947) );
  AN2 C6265 ( .A(n1945), .B(n1492), .Z(n1946) );
  AN2 C6266 ( .A(n1944), .B(n1554), .Z(n1945) );
  AN2 C6267 ( .A(n1943), .B(n1610), .Z(n1944) );
  AN2 C6268 ( .A(n1942), .B(n1720), .Z(n1943) );
  AN2 C6269 ( .A(n1941), .B(n1660), .Z(n1942) );
  AN2 C6270 ( .A(n1940), .B(n1783), .Z(n1941) );
  AN2 C6271 ( .A(n1939), .B(n1815), .Z(n1940) );
  AN2 C6272 ( .A(n1938), .B(n1857), .Z(n1939) );
  AN2 C6273 ( .A(n1937), .B(n1850), .Z(n1938) );
  AN2 C6274 ( .A(n1846), .B(n1268), .Z(n1937) );
  AN2 C6276 ( .A(n1955), .B(n1308), .Z(n119) );
  AN2 C6277 ( .A(n1954), .B(n1410), .Z(n1955) );
  AN2 C6278 ( .A(n1953), .B(n1480), .Z(n1954) );
  AN2 C6279 ( .A(n1952), .B(n1540), .Z(n1953) );
  AN2 C6280 ( .A(n1951), .B(n1596), .Z(n1952) );
  AN2 C6281 ( .A(n1950), .B(n1704), .Z(n1951) );
  AN2 C6282 ( .A(n1949), .B(n1648), .Z(n1950) );
  AN2 C6283 ( .A(n1948), .B(n1768), .Z(n1949) );
  AN2 C6284 ( .A(n1843), .B(n1809), .Z(n1948) );
  AN2 C6286 ( .A(n1963), .B(n1288), .Z(n120) );
  AN2 C6287 ( .A(n1962), .B(n1384), .Z(n1963) );
  AN2 C6288 ( .A(n1961), .B(n1468), .Z(n1962) );
  AN2 C6289 ( .A(n1960), .B(n1526), .Z(n1961) );
  AN2 C6290 ( .A(n1959), .B(n1582), .Z(n1960) );
  AN2 C62911 ( .A(n1958), .B(n1688), .Z(n1959) );
  AN2 C6292 ( .A(n1957), .B(n1636), .Z(n1958) );
  AN2 C6293 ( .A(n1956), .B(n1752), .Z(n1957) );
  AN2 C6294 ( .A(n1840), .B(n1803), .Z(n1956) );
  AN2 C6296 ( .A(n1971), .B(n1278), .Z(n121) );
  AN2 C6297 ( .A(n1970), .B(n1371), .Z(n1971) );
  AN2 C6298 ( .A(n1969), .B(n1462), .Z(n1970) );
  AN2 C6299 ( .A(n1968), .B(n1519), .Z(n1969) );
  AN2 C6300 ( .A(n1967), .B(n1575), .Z(n1968) );
  AN2 C6301 ( .A(n1966), .B(n1680), .Z(n1967) );
  AN2 C6302 ( .A(n1965), .B(n1630), .Z(n1966) );
  AN2 C6303 ( .A(n1964), .B(n1744), .Z(n1965) );
  AN2 C6304 ( .A(n1837), .B(n1800), .Z(n1964) );
  AN2 C6306 ( .A(n1982), .B(n1358), .Z(n122) );
  AN2 C6307 ( .A(n1981), .B(n1456), .Z(n1982) );
  AN2 C6308 ( .A(n1980), .B(n1512), .Z(n1981) );
  AN2 C6309 ( .A(n1979), .B(n1568), .Z(n1980) );
  AN2 C6310 ( .A(n1978), .B(n1624), .Z(n1979) );
  AN2 C63111 ( .A(n1977), .B(n1736), .Z(n1978) );
  AN2 C63121 ( .A(n1976), .B(n1672), .Z(n1977) );
  AN2 C6313 ( .A(n1975), .B(n1798), .Z(n1976) );
  AN2 C6314 ( .A(n1974), .B(n1821), .Z(n1975) );
  AN2 C6315 ( .A(n1973), .B(n1868), .Z(n1974) );
  AN2 C6316 ( .A(n1972), .B(n1861), .Z(n1973) );
  AN2 C6317 ( .A(n1834), .B(n1349), .Z(n1972) );
  AN2 C6319 ( .A(n1990), .B(n1337), .Z(n123) );
  AN2 C6320 ( .A(n1989), .B(n1446), .Z(n1990) );
  AN2 C63211 ( .A(n1988), .B(n1498), .Z(n1989) );
  AN2 C63221 ( .A(n1987), .B(n1561), .Z(n1988) );
  AN2 C6323 ( .A(n1986), .B(n1617), .Z(n1987) );
  AN2 C6324 ( .A(n1985), .B(n1728), .Z(n1986) );
  AN2 C6325 ( .A(n1984), .B(n1666), .Z(n1985) );
  AN2 C6326 ( .A(n1983), .B(n1791), .Z(n1984) );
  AN2 C6327 ( .A(n1831), .B(n1818), .Z(n1983) );
  AN2 C6329 ( .A(n1998), .B(n1318), .Z(n124) );
  AN2 C6330 ( .A(n1997), .B(n1423), .Z(n1998) );
  AN2 C6331 ( .A(n1996), .B(n1486), .Z(n1997) );
  AN2 C6332 ( .A(n1995), .B(n1547), .Z(n1996) );
  AN2 C6333 ( .A(n1994), .B(n1603), .Z(n1995) );
  AN2 C6334 ( .A(n1993), .B(n1712), .Z(n1994) );
  AN2 C6335 ( .A(n1992), .B(n1654), .Z(n1993) );
  AN2 C6336 ( .A(n1991), .B(n1776), .Z(n1992) );
  AN2 C6337 ( .A(n1828), .B(n1812), .Z(n1991) );
  AN2 C6339 ( .A(n2006), .B(n1298), .Z(n125) );
  AN2 C6340 ( .A(n2005), .B(n1397), .Z(n2006) );
  AN2 C63411 ( .A(n2004), .B(n1474), .Z(n2005) );
  AN2 C6342 ( .A(n2003), .B(n1533), .Z(n2004) );
  AN2 C6343 ( .A(n2002), .B(n1589), .Z(n2003) );
  AN2 C6344 ( .A(n2001), .B(n1696), .Z(n2002) );
  AN2 C6345 ( .A(n2000), .B(n1642), .Z(n2001) );
  AN2 C6346 ( .A(n1999), .B(n1760), .Z(n2000) );
  AN2 C6347 ( .A(n1825), .B(n1806), .Z(n1999) );
  OR2 C6349 ( .A(n2019), .B(n2020), .Z(n126) );
  OR2 C6350 ( .A(n2017), .B(n2018), .Z(n2019) );
  OR2 C6351 ( .A(n2015), .B(n2016), .Z(n2017) );
  OR2 C6352 ( .A(n2013), .B(n2014), .Z(n2015) );
  OR2 C6353 ( .A(n2011), .B(n2012), .Z(n2013) );
  OR2 C6354 ( .A(n2009), .B(n2010), .Z(n2011) );
  OR2 C6355 ( .A(n2007), .B(n2008), .Z(n2009) );
  AN2 C6356 ( .A(n125), .B(U154_Z_5), .Z(n2007) );
  AN2 C6357 ( .A(n124), .B(U154_Z_4), .Z(n2008) );
  AN2 C6358 ( .A(n123), .B(U154_Z_3), .Z(n2010) );
  AN2 C6359 ( .A(n122), .B(U155_Z_1), .Z(n2012) );
  AN2 C6360 ( .A(n121), .B(U154_Z_2), .Z(n2014) );
  AN2 C63611 ( .A(n120), .B(U154_Z_1), .Z(n2016) );
  AN2 C6362 ( .A(n119), .B(U154_Z_0), .Z(n2018) );
  AN2 C6363 ( .A(n110), .B(U155_Z_0), .Z(n2020) );
  AN2 C6724 ( .A(U155_Z_0), .B(n5303), .Z(n255) );
  AN2 C6726 ( .A(U154_Z_0), .B(n5323), .Z(n257) );
  AN2 C6728 ( .A(U154_Z_1), .B(n5341), .Z(n259) );
  AN2 C6730 ( .A(U154_Z_2), .B(n5359), .Z(n261) );
  AN2 C6732 ( .A(U155_Z_1), .B(n5378), .Z(n263) );
  AN2 C6734 ( .A(U154_Z_3), .B(n5398), .Z(n265) );
  AN2 C6736 ( .A(U154_Z_4), .B(n5416), .Z(n267) );
  AN2 C6738 ( .A(U154_Z_5), .B(n5434), .Z(n269) );
  AN2 C6740 ( .A(U155_Z_0), .B(n2021), .Z(n271) );
  OR2 C6741 ( .A(n5307), .B(n5315), .Z(n2021) );
  AN2 C6743 ( .A(U155_Z_0), .B(n5315), .Z(n273) );
  AN2 C6745 ( .A(U155_Z_1), .B(n2022), .Z(n275) );
  OR2 C6746 ( .A(n5382), .B(n5390), .Z(n2022) );
  AN2 C6748 ( .A(U155_Z_1), .B(n5390), .Z(n277) );
  AN2 C6750 ( .A(U155_Z_0), .B(n5302), .Z(n279) );
  AN2 C6752 ( .A(U155_Z_1), .B(n5377), .Z(n281) );
  AN2 C6754 ( .A(U155_Z_0), .B(n2030), .Z(n283) );
  OR2 C6755 ( .A(n2029), .B(n5314), .Z(n2030) );
  OR2 C6756 ( .A(n2028), .B(n5313), .Z(n2029) );
  OR2 C6757 ( .A(n2027), .B(n5305), .Z(n2028) );
  OR2 C6758 ( .A(n2026), .B(n5312), .Z(n2027) );
  OR2 C6759 ( .A(n2025), .B(n5311), .Z(n2026) );
  OR2 C6760 ( .A(n2024), .B(n5309), .Z(n2025) );
  OR2 C6761 ( .A(n2023), .B(n5310), .Z(n2024) );
  OR2 C6762 ( .A(n5304), .B(n5308), .Z(n2023) );
  AN2 C6764 ( .A(U154_Z_0), .B(n2038), .Z(n285) );
  OR2 C6765 ( .A(n2037), .B(n5333), .Z(n2038) );
  OR2 C6766 ( .A(n2036), .B(n5332), .Z(n2037) );
  OR2 C6767 ( .A(n2035), .B(n5325), .Z(n2036) );
  OR2 C6768 ( .A(n2034), .B(n5331), .Z(n2035) );
  OR2 C6769 ( .A(n2033), .B(n5330), .Z(n2034) );
  OR2 C6770 ( .A(n2032), .B(n5328), .Z(n2033) );
  OR2 C67711 ( .A(n2031), .B(n5329), .Z(n2032) );
  OR2 C6772 ( .A(n5324), .B(n5327), .Z(n2031) );
  AN2 C6774 ( .A(U154_Z_1), .B(n2046), .Z(n287) );
  OR2 C6775 ( .A(n2045), .B(n5351), .Z(n2046) );
  OR2 C6776 ( .A(n2044), .B(n5350), .Z(n2045) );
  OR2 C6777 ( .A(n2043), .B(n5343), .Z(n2044) );
  OR2 C6778 ( .A(n2042), .B(n5349), .Z(n2043) );
  OR2 C6779 ( .A(n2041), .B(n5348), .Z(n2042) );
  OR2 C6780 ( .A(n2040), .B(n5346), .Z(n2041) );
  OR2 C67811 ( .A(n2039), .B(n5347), .Z(n2040) );
  OR2 C6782 ( .A(n5342), .B(n5345), .Z(n2039) );
  AN2 C6784 ( .A(U154_Z_2), .B(n2054), .Z(n289) );
  OR2 C6785 ( .A(n2053), .B(n5369), .Z(n2054) );
  OR2 C6786 ( .A(n2052), .B(n5368), .Z(n2053) );
  OR2 C6787 ( .A(n2051), .B(n5361), .Z(n2052) );
  OR2 C6788 ( .A(n2050), .B(n5367), .Z(n2051) );
  OR2 C6789 ( .A(n2049), .B(n5366), .Z(n2050) );
  OR2 C6790 ( .A(n2048), .B(n5364), .Z(n2049) );
  OR2 C67911 ( .A(n2047), .B(n5365), .Z(n2048) );
  OR2 C6792 ( .A(n5360), .B(n5363), .Z(n2047) );
  AN2 C6794 ( .A(U155_Z_1), .B(n2062), .Z(n291) );
  OR2 C6795 ( .A(n2061), .B(n5389), .Z(n2062) );
  OR2 C6796 ( .A(n2060), .B(n5388), .Z(n2061) );
  OR2 C6797 ( .A(n2059), .B(n5380), .Z(n2060) );
  OR2 C6798 ( .A(n2058), .B(n5387), .Z(n2059) );
  OR2 C6799 ( .A(n2057), .B(n5386), .Z(n2058) );
  OR2 C6800 ( .A(n2056), .B(n5384), .Z(n2057) );
  OR2 C68011 ( .A(n2055), .B(n5385), .Z(n2056) );
  OR2 C6802 ( .A(n5379), .B(n5383), .Z(n2055) );
  AN2 C6804 ( .A(U154_Z_3), .B(n2070), .Z(n293) );
  OR2 C6805 ( .A(n2069), .B(n5408), .Z(n2070) );
  OR2 C6806 ( .A(n2068), .B(n5407), .Z(n2069) );
  OR2 C6807 ( .A(n2067), .B(n5400), .Z(n2068) );
  OR2 C6808 ( .A(n2066), .B(n5406), .Z(n2067) );
  OR2 C6809 ( .A(n2065), .B(n5405), .Z(n2066) );
  OR2 C6810 ( .A(n2064), .B(n5403), .Z(n2065) );
  OR2 C68111 ( .A(n2063), .B(n5404), .Z(n2064) );
  OR2 C6812 ( .A(n5399), .B(n5402), .Z(n2063) );
  AN2 C6814 ( .A(U154_Z_4), .B(n2078), .Z(n295) );
  OR2 C6815 ( .A(n2077), .B(n5426), .Z(n2078) );
  OR2 C6816 ( .A(n2076), .B(n5425), .Z(n2077) );
  OR2 C6817 ( .A(n2075), .B(n5418), .Z(n2076) );
  OR2 C6818 ( .A(n2074), .B(n5424), .Z(n2075) );
  OR2 C6819 ( .A(n2073), .B(n5423), .Z(n2074) );
  OR2 C6820 ( .A(n2072), .B(n5421), .Z(n2073) );
  OR2 C68211 ( .A(n2071), .B(n5422), .Z(n2072) );
  OR2 C6822 ( .A(n5417), .B(n5420), .Z(n2071) );
  AN2 C6824 ( .A(U154_Z_5), .B(n2086), .Z(n297) );
  OR2 C6825 ( .A(n2085), .B(n5444), .Z(n2086) );
  OR2 C6826 ( .A(n2084), .B(n5443), .Z(n2085) );
  OR2 C6827 ( .A(n2083), .B(n5436), .Z(n2084) );
  OR2 C6828 ( .A(n2082), .B(n5442), .Z(n2083) );
  OR2 C6829 ( .A(n2081), .B(n5441), .Z(n2082) );
  OR2 C6830 ( .A(n2080), .B(n5439), .Z(n2081) );
  OR2 C68311 ( .A(n2079), .B(n5440), .Z(n2080) );
  OR2 C6832 ( .A(n5435), .B(n5438), .Z(n2079) );
  AN2 C6834 ( .A(n2088), .B(n289), .Z(n299) );
  AN2 C6835 ( .A(n2087), .B(n287), .Z(n2088) );
  AN2 C6836 ( .A(n283), .B(n285), .Z(n2087) );
  AN2 C6837 ( .A(n2090), .B(n5297), .Z(n300) );
  AN2 C6838 ( .A(n2089), .B(n5296), .Z(n2090) );
  AN2 C6839 ( .A(n271), .B(n5295), .Z(n2089) );
  AN2 C6840 ( .A(n5274), .B(n5295), .Z(n301) );
  AN2 C6841 ( .A(n301), .B(n5296), .Z(n302) );
  AN2 C6842 ( .A(n302), .B(n261), .Z(n303) );
  AN2 C6843 ( .A(n302), .B(n5297), .Z(n304) );
  AN2 C6844 ( .A(n304), .B(n5298), .Z(n305) );
  AN2 C6845 ( .A(n305), .B(n5299), .Z(n306) );
  AN2 C6846 ( .A(n2093), .B(n297), .Z(n307) );
  AN2 C6847 ( .A(n2092), .B(n295), .Z(n2093) );
  AN2 C6848 ( .A(n2091), .B(n293), .Z(n2092) );
  AN2 C6849 ( .A(n299), .B(n291), .Z(n2091) );
  AN2 C6850 ( .A(n2096), .B(n5301), .Z(n308) );
  AN2 C6851 ( .A(n2095), .B(n5300), .Z(n2096) );
  AN2 C6852 ( .A(n2094), .B(n5299), .Z(n2095) );
  AN2 C6853 ( .A(n299), .B(n275), .Z(n2094) );
  AN2 C6854 ( .A(n2099), .B(n5301), .Z(n309) );
  AN2 C6855 ( .A(n2098), .B(n5300), .Z(n2099) );
  AN2 C6856 ( .A(n2097), .B(n5299), .Z(n2098) );
  AN2 C6857 ( .A(n299), .B(n281), .Z(n2097) );
  AN2 C6858 ( .A(n2102), .B(n5301), .Z(n310) );
  AN2 C6859 ( .A(n2101), .B(n5300), .Z(n2102) );
  AN2 C6860 ( .A(n2100), .B(n5299), .Z(n2101) );
  AN2 C6861 ( .A(n300), .B(n281), .Z(n2100) );
  AN2 C6862 ( .A(n2105), .B(n5301), .Z(n311) );
  AN2 C6863 ( .A(n2104), .B(n5300), .Z(n2105) );
  AN2 C6864 ( .A(n2103), .B(n5299), .Z(n2104) );
  AN2 C6865 ( .A(n300), .B(n275), .Z(n2103) );
  AN2 C6866 ( .A(n2111), .B(n5301), .Z(n312) );
  AN2 C6867 ( .A(n2110), .B(n5300), .Z(n2111) );
  AN2 C6868 ( .A(n2109), .B(n5299), .Z(n2110) );
  AN2 C6869 ( .A(n2108), .B(n5298), .Z(n2109) );
  AN2 C6870 ( .A(n2107), .B(n5297), .Z(n2108) );
  AN2 C68711 ( .A(n2106), .B(n5296), .Z(n2107) );
  AN2 C6872 ( .A(n279), .B(n5295), .Z(n2106) );
  AN2 C6873 ( .A(n2114), .B(n297), .Z(n313) );
  AN2 C6874 ( .A(n2113), .B(n295), .Z(n2114) );
  AN2 C6875 ( .A(n2112), .B(n293), .Z(n2113) );
  AN2 C6876 ( .A(n300), .B(n291), .Z(n2112) );
  AN2 C6877 ( .A(n2120), .B(n297), .Z(n314) );
  AN2 C6878 ( .A(n2119), .B(n295), .Z(n2120) );
  AN2 C6879 ( .A(n2118), .B(n293), .Z(n2119) );
  AN2 C6880 ( .A(n2117), .B(n291), .Z(n2118) );
  AN2 C68811 ( .A(n2116), .B(n289), .Z(n2117) );
  AN2 C6882 ( .A(n2115), .B(n287), .Z(n2116) );
  AN2 C6883 ( .A(n255), .B(n285), .Z(n2115) );
  AN2 C6884 ( .A(n2126), .B(n297), .Z(n315) );
  AN2 C6885 ( .A(n2125), .B(n295), .Z(n2126) );
  AN2 C6886 ( .A(n2124), .B(n293), .Z(n2125) );
  AN2 C6887 ( .A(n2123), .B(n291), .Z(n2124) );
  AN2 C6888 ( .A(n2122), .B(n289), .Z(n2123) );
  AN2 C6889 ( .A(n2121), .B(n287), .Z(n2122) );
  AN2 C6890 ( .A(n5274), .B(n257), .Z(n2121) );
  AN2 C68911 ( .A(n2131), .B(n297), .Z(n316) );
  AN2 C6892 ( .A(n2130), .B(n295), .Z(n2131) );
  AN2 C6893 ( .A(n2129), .B(n293), .Z(n2130) );
  AN2 C6894 ( .A(n2128), .B(n291), .Z(n2129) );
  AN2 C6895 ( .A(n2127), .B(n289), .Z(n2128) );
  AN2 C6896 ( .A(n301), .B(n259), .Z(n2127) );
  AN2 C6897 ( .A(n2135), .B(n2136), .Z(n317) );
  AN2 C6898 ( .A(n2134), .B(n297), .Z(n2135) );
  AN2 C6899 ( .A(n2133), .B(n295), .Z(n2134) );
  AN2 C6900 ( .A(n2132), .B(n293), .Z(n2133) );
  AN2 C69011 ( .A(n303), .B(n291), .Z(n2132) );
  IV I_1861 ( .A(ALTERNATE_ENCODE), .Z(n2136) );
  AN2 C6903 ( .A(n2140), .B(ALTERNATE_ENCODE), .Z(n318) );
  AN2 C6904 ( .A(n2139), .B(n5301), .Z(n2140) );
  AN2 C6905 ( .A(n2138), .B(n5300), .Z(n2139) );
  AN2 C6906 ( .A(n2137), .B(n5299), .Z(n2138) );
  AN2 C6907 ( .A(n303), .B(n275), .Z(n2137) );
  AN2 C6908 ( .A(n2143), .B(n297), .Z(n319) );
  AN2 C6909 ( .A(n2142), .B(n295), .Z(n2143) );
  AN2 C6910 ( .A(n2141), .B(n293), .Z(n2142) );
  AN2 C69111 ( .A(n304), .B(n263), .Z(n2141) );
  AN2 C6912 ( .A(n2145), .B(n297), .Z(n320) );
  AN2 C6913 ( .A(n2144), .B(n295), .Z(n2145) );
  AN2 C6914 ( .A(n305), .B(n265), .Z(n2144) );
  AN2 C6915 ( .A(n2146), .B(n297), .Z(n321) );
  AN2 C6916 ( .A(n306), .B(n267), .Z(n2146) );
  AN2 C6917 ( .A(n2147), .B(n269), .Z(n322) );
  AN2 C6918 ( .A(n306), .B(n5300), .Z(n2147) );
  AN2 C7050 ( .A(n97), .B(n5627), .Z(n749) );
  IV I_239 ( .A(test_pat_seed_a[57]), .Z(U37_DATA4_57) );
  IV I_240 ( .A(test_pat_seed_a[56]), .Z(U37_DATA4_56) );
  IV I_2411 ( .A(test_pat_seed_a[55]), .Z(U37_DATA4_55) );
  IV I_2421 ( .A(test_pat_seed_a[54]), .Z(U37_DATA4_54) );
  IV I_2431 ( .A(test_pat_seed_a[53]), .Z(U37_DATA4_53) );
  IV I_244 ( .A(test_pat_seed_a[52]), .Z(U37_DATA4_52) );
  IV I_245 ( .A(test_pat_seed_a[51]), .Z(U37_DATA4_51) );
  IV I_246 ( .A(test_pat_seed_a[50]), .Z(U37_DATA4_50) );
  IV I_247 ( .A(test_pat_seed_a[49]), .Z(U37_DATA4_49) );
  IV I_248 ( .A(test_pat_seed_a[48]), .Z(U37_DATA4_48) );
  IV I_249 ( .A(test_pat_seed_a[47]), .Z(U37_DATA4_47) );
  IV I_250 ( .A(test_pat_seed_a[46]), .Z(U37_DATA4_46) );
  IV I_2511 ( .A(test_pat_seed_a[45]), .Z(U37_DATA4_45) );
  IV I_2521 ( .A(test_pat_seed_a[44]), .Z(U37_DATA4_44) );
  IV I_2531 ( .A(test_pat_seed_a[43]), .Z(U37_DATA4_43) );
  IV I_254 ( .A(test_pat_seed_a[42]), .Z(U37_DATA4_42) );
  IV I_255 ( .A(test_pat_seed_a[41]), .Z(U37_DATA4_41) );
  IV I_256 ( .A(test_pat_seed_a[40]), .Z(U37_DATA4_40) );
  IV I_257 ( .A(test_pat_seed_a[39]), .Z(U37_DATA4_39) );
  IV I_258 ( .A(test_pat_seed_a[38]), .Z(U37_DATA4_38) );
  IV I_259 ( .A(test_pat_seed_a[37]), .Z(U37_DATA4_37) );
  IV I_260 ( .A(test_pat_seed_a[36]), .Z(U37_DATA4_36) );
  IV I_2611 ( .A(test_pat_seed_a[35]), .Z(U37_DATA4_35) );
  IV I_2621 ( .A(test_pat_seed_a[34]), .Z(U37_DATA4_34) );
  IV I_2631 ( .A(test_pat_seed_a[33]), .Z(U37_DATA4_33) );
  IV I_264 ( .A(test_pat_seed_a[32]), .Z(U37_DATA4_32) );
  IV I_265 ( .A(test_pat_seed_a[31]), .Z(U37_DATA4_31) );
  IV I_266 ( .A(test_pat_seed_a[30]), .Z(U37_DATA4_30) );
  IV I_267 ( .A(test_pat_seed_a[29]), .Z(U37_DATA4_29) );
  IV I_268 ( .A(test_pat_seed_a[28]), .Z(U37_DATA4_28) );
  IV I_269 ( .A(test_pat_seed_a[27]), .Z(U37_DATA4_27) );
  IV I_270 ( .A(test_pat_seed_a[26]), .Z(U37_DATA4_26) );
  IV I_2711 ( .A(test_pat_seed_a[25]), .Z(U37_DATA4_25) );
  IV I_2721 ( .A(test_pat_seed_a[24]), .Z(U37_DATA4_24) );
  IV I_2731 ( .A(test_pat_seed_a[23]), .Z(U37_DATA4_23) );
  IV I_274 ( .A(test_pat_seed_a[22]), .Z(U37_DATA4_22) );
  IV I_275 ( .A(test_pat_seed_a[21]), .Z(U37_DATA4_21) );
  IV I_276 ( .A(test_pat_seed_a[20]), .Z(U37_DATA4_20) );
  IV I_277 ( .A(test_pat_seed_a[19]), .Z(U37_DATA4_19) );
  IV I_278 ( .A(test_pat_seed_a[18]), .Z(U37_DATA4_18) );
  IV I_279 ( .A(test_pat_seed_a[17]), .Z(U37_DATA4_17) );
  IV I_280 ( .A(test_pat_seed_a[16]), .Z(U37_DATA4_16) );
  IV I_2811 ( .A(test_pat_seed_a[15]), .Z(U37_DATA4_15) );
  IV I_2821 ( .A(test_pat_seed_a[14]), .Z(U37_DATA4_14) );
  IV I_2831 ( .A(test_pat_seed_a[13]), .Z(U37_DATA4_13) );
  IV I_284 ( .A(test_pat_seed_a[12]), .Z(U37_DATA4_12) );
  IV I_285 ( .A(test_pat_seed_a[11]), .Z(U37_DATA4_11) );
  IV I_286 ( .A(test_pat_seed_a[10]), .Z(U37_DATA4_10) );
  IV I_287 ( .A(test_pat_seed_a[9]), .Z(U37_DATA4_9) );
  IV I_288 ( .A(test_pat_seed_a[8]), .Z(U37_DATA4_8) );
  IV I_289 ( .A(test_pat_seed_a[7]), .Z(U37_DATA4_7) );
  IV I_290 ( .A(test_pat_seed_a[6]), .Z(U37_DATA4_6) );
  IV I_2911 ( .A(test_pat_seed_a[5]), .Z(U37_DATA4_5) );
  IV I_2921 ( .A(test_pat_seed_a[4]), .Z(U37_DATA4_4) );
  IV I_293 ( .A(test_pat_seed_a[3]), .Z(U37_DATA4_3) );
  IV I_294 ( .A(test_pat_seed_a[2]), .Z(U37_DATA4_2) );
  IV I_295 ( .A(test_pat_seed_a[1]), .Z(U37_DATA4_1) );
  IV I_296 ( .A(test_pat_seed_a[0]), .Z(U37_DATA4_0) );
  IV I_297 ( .A(test_pat_seed_b[57]), .Z(U37_DATA6_57) );
  IV I_298 ( .A(test_pat_seed_b[56]), .Z(U37_DATA6_56) );
  IV I_299 ( .A(test_pat_seed_b[55]), .Z(U37_DATA6_55) );
  IV I_300 ( .A(test_pat_seed_b[54]), .Z(U37_DATA6_54) );
  IV I_3011 ( .A(test_pat_seed_b[53]), .Z(U37_DATA6_53) );
  IV I_3021 ( .A(test_pat_seed_b[52]), .Z(U37_DATA6_52) );
  IV I_303 ( .A(test_pat_seed_b[51]), .Z(U37_DATA6_51) );
  IV I_304 ( .A(test_pat_seed_b[50]), .Z(U37_DATA6_50) );
  IV I_305 ( .A(test_pat_seed_b[49]), .Z(U37_DATA6_49) );
  IV I_306 ( .A(test_pat_seed_b[48]), .Z(U37_DATA6_48) );
  IV I_307 ( .A(test_pat_seed_b[47]), .Z(U37_DATA6_47) );
  IV I_308 ( .A(test_pat_seed_b[46]), .Z(U37_DATA6_46) );
  IV I_309 ( .A(test_pat_seed_b[45]), .Z(U37_DATA6_45) );
  IV I_3101 ( .A(test_pat_seed_b[44]), .Z(U37_DATA6_44) );
  IV I_3111 ( .A(test_pat_seed_b[43]), .Z(U37_DATA6_43) );
  IV I_3121 ( .A(test_pat_seed_b[42]), .Z(U37_DATA6_42) );
  IV I_3131 ( .A(test_pat_seed_b[41]), .Z(U37_DATA6_41) );
  IV I_3141 ( .A(test_pat_seed_b[40]), .Z(U37_DATA6_40) );
  IV I_3151 ( .A(test_pat_seed_b[39]), .Z(U37_DATA6_39) );
  IV I_316 ( .A(test_pat_seed_b[38]), .Z(U37_DATA6_38) );
  IV I_317 ( .A(test_pat_seed_b[37]), .Z(U37_DATA6_37) );
  IV I_318 ( .A(test_pat_seed_b[36]), .Z(U37_DATA6_36) );
  IV I_319 ( .A(test_pat_seed_b[35]), .Z(U37_DATA6_35) );
  IV I_320 ( .A(test_pat_seed_b[34]), .Z(U37_DATA6_34) );
  IV I_3211 ( .A(test_pat_seed_b[33]), .Z(U37_DATA6_33) );
  IV I_3221 ( .A(test_pat_seed_b[32]), .Z(U37_DATA6_32) );
  IV I_323 ( .A(test_pat_seed_b[31]), .Z(U37_DATA6_31) );
  IV I_324 ( .A(test_pat_seed_b[30]), .Z(U37_DATA6_30) );
  IV I_325 ( .A(test_pat_seed_b[29]), .Z(U37_DATA6_29) );
  IV I_326 ( .A(test_pat_seed_b[28]), .Z(U37_DATA6_28) );
  IV I_327 ( .A(test_pat_seed_b[27]), .Z(U37_DATA6_27) );
  IV I_328 ( .A(test_pat_seed_b[26]), .Z(U37_DATA6_26) );
  IV I_329 ( .A(test_pat_seed_b[25]), .Z(U37_DATA6_25) );
  IV I_330 ( .A(test_pat_seed_b[24]), .Z(U37_DATA6_24) );
  IV I_3311 ( .A(test_pat_seed_b[23]), .Z(U37_DATA6_23) );
  IV I_3321 ( .A(test_pat_seed_b[22]), .Z(U37_DATA6_22) );
  IV I_333 ( .A(test_pat_seed_b[21]), .Z(U37_DATA6_21) );
  IV I_334 ( .A(test_pat_seed_b[20]), .Z(U37_DATA6_20) );
  IV I_335 ( .A(test_pat_seed_b[19]), .Z(U37_DATA6_19) );
  IV I_336 ( .A(test_pat_seed_b[18]), .Z(U37_DATA6_18) );
  IV I_337 ( .A(test_pat_seed_b[17]), .Z(U37_DATA6_17) );
  IV I_338 ( .A(test_pat_seed_b[16]), .Z(U37_DATA6_16) );
  IV I_339 ( .A(test_pat_seed_b[15]), .Z(U37_DATA6_15) );
  IV I_340 ( .A(test_pat_seed_b[14]), .Z(U37_DATA6_14) );
  IV I_3411 ( .A(test_pat_seed_b[13]), .Z(U37_DATA6_13) );
  IV I_3421 ( .A(test_pat_seed_b[12]), .Z(U37_DATA6_12) );
  IV I_343 ( .A(test_pat_seed_b[11]), .Z(U37_DATA6_11) );
  IV I_344 ( .A(test_pat_seed_b[10]), .Z(U37_DATA6_10) );
  IV I_345 ( .A(test_pat_seed_b[9]), .Z(U37_DATA6_9) );
  IV I_346 ( .A(test_pat_seed_b[8]), .Z(U37_DATA6_8) );
  IV I_347 ( .A(test_pat_seed_b[7]), .Z(U37_DATA6_7) );
  IV I_348 ( .A(test_pat_seed_b[6]), .Z(U37_DATA6_6) );
  IV I_349 ( .A(test_pat_seed_b[5]), .Z(U37_DATA6_5) );
  IV I_350 ( .A(test_pat_seed_b[4]), .Z(U37_DATA6_4) );
  IV I_3511 ( .A(test_pat_seed_b[3]), .Z(U37_DATA6_3) );
  IV I_3521 ( .A(test_pat_seed_b[2]), .Z(U37_DATA6_2) );
  IV I_353 ( .A(test_pat_seed_b[1]), .Z(U37_DATA6_1) );
  IV I_354 ( .A(test_pat_seed_b[0]), .Z(U37_DATA6_0) );
  IV I_356 ( .A(reset_to_pma_tx), .Z(n1148) );
  AN2 C198 ( .A(n5527), .B(n5526), .Z(n2533) );
  AN2 C19910 ( .A(n5525), .B(n5517), .Z(n2534) );
  OR2 C203 ( .A(n5527), .B(U112_DATA3_0), .Z(n2536) );
  OR2 C2043 ( .A(U113_DATA3_0), .B(n5517), .Z(n2537) );
  OR2 C2091 ( .A(U111_DATA3_0), .B(n5526), .Z(n2540) );
  OR2 C2101 ( .A(n5525), .B(U114_DATA2_0), .Z(n2541) );
  OR2 C2151 ( .A(n5527), .B(U112_DATA3_0), .Z(n2544) );
  OR2 C2161 ( .A(n5525), .B(U114_DATA2_0), .Z(n2545) );
  AN2 C2191 ( .A(U111_DATA3_0), .B(U112_DATA3_0), .Z(n2548) );
  AN2 C220 ( .A(U113_DATA3_0), .B(U114_DATA2_0), .Z(n2549) );
  OR2 C224 ( .A(U111_DATA3_0), .B(U112_DATA3_0), .Z(n2551) );
  OR2 C225 ( .A(n5525), .B(n5517), .Z(n2552) );
  OR2 C230 ( .A(n5527), .B(n5526), .Z(n2555) );
  OR2 C231 ( .A(U113_DATA3_0), .B(U114_DATA2_0), .Z(n2556) );
  OR2 C236 ( .A(U111_DATA3_0), .B(n5526), .Z(n2559) );
  OR2 C237 ( .A(U113_DATA3_0), .B(n5517), .Z(n2560) );
  OR2 C243 ( .A(U111_DATA3_0), .B(n5526), .Z(n2563) );
  OR2 C244 ( .A(n5525), .B(n5517), .Z(n2564) );
  OR2 C249 ( .A(n5527), .B(U112_DATA3_0), .Z(n2566) );
  OR2 C250 ( .A(n5525), .B(n5517), .Z(n2567) );
  OR2 C255 ( .A(n5527), .B(n5526), .Z(n2569) );
  OR2 C256 ( .A(U113_DATA3_0), .B(n5517), .Z(n2570) );
  OR2 C259 ( .A(U111_DATA3_0), .B(U112_DATA3_0), .Z(n2572) );
  OR2 C260 ( .A(U113_DATA3_0), .B(n5517), .Z(n2573) );
  OR2 C265 ( .A(n5527), .B(n5526), .Z(n2575) );
  OR2 C266 ( .A(n5525), .B(U114_DATA2_0), .Z(n2576) );
  OR2 C269 ( .A(U111_DATA3_0), .B(U112_DATA3_0), .Z(n2578) );
  OR2 C2701 ( .A(n5525), .B(U114_DATA2_0), .Z(n2579) );
  OR2 C273 ( .A(U111_DATA3_0), .B(n5526), .Z(n2581) );
  OR2 C274 ( .A(U113_DATA3_0), .B(U114_DATA2_0), .Z(n2582) );
  OR2 C277 ( .A(n5527), .B(U112_DATA3_0), .Z(n2584) );
  OR2 C278 ( .A(U113_DATA3_0), .B(U114_DATA2_0), .Z(n2585) );
  AN2 C4802 ( .A(U3_U1_DATA1_14), .B(U3_U1_DATA1_15), .Z(n2675) );
  AN2 C4811 ( .A(U3_U1_DATA1_13), .B(n2675), .Z(n2676) );
  AN2 C4821 ( .A(U3_U1_DATA1_12), .B(n2676), .Z(n2677) );
  AN2 C483 ( .A(U3_U1_DATA1_11), .B(n2677), .Z(n2678) );
  AN2 C4841 ( .A(U3_U1_DATA1_10), .B(n2678), .Z(n2679) );
  AN2 C485 ( .A(U3_U1_DATA1_9), .B(n2679), .Z(n2680) );
  AN2 C4861 ( .A(U3_U1_DATA1_8), .B(n2680), .Z(n2681) );
  AN2 C4871 ( .A(U3_U1_DATA1_7), .B(n2681), .Z(n2682) );
  AN2 C488 ( .A(U3_U1_DATA1_6), .B(n2682), .Z(n2683) );
  AN2 C489 ( .A(U3_U1_DATA1_5), .B(n2683), .Z(n2684) );
  AN2 C490 ( .A(U3_U1_DATA1_4), .B(n2684), .Z(n2685) );
  AN2 C4911 ( .A(U3_U1_DATA1_3), .B(n2685), .Z(n2686) );
  AN2 C4921 ( .A(U3_U1_DATA1_2), .B(n2686), .Z(n2687) );
  AN2 C4932 ( .A(U3_U1_DATA1_1), .B(n2687), .Z(n2688) );
  AN2 C4941 ( .A(U3_U1_DATA1_0), .B(n2688), .Z(n2689) );
  OR2 C4952 ( .A(sub_128_aco_A_7_), .B(sub_128_aco_A_8_), .Z(n2690) );
  OR2 C4961 ( .A(sub_128_aco_A_6_), .B(n2690), .Z(n2691) );
  OR2 C4972 ( .A(sub_128_aco_A_5_), .B(n2691), .Z(n2692) );
  OR2 C498 ( .A(sub_128_aco_A_4_), .B(n2692), .Z(n2693) );
  OR2 C4991 ( .A(sub_128_aco_A_3_), .B(n2693), .Z(n2694) );
  OR2 C500 ( .A(sub_128_aco_A_2_), .B(n2694), .Z(n2695) );
  OR2 C5011 ( .A(sub_128_aco_A_1_), .B(n2695), .Z(n2696) );
  OR2 C502 ( .A(sub_128_aco_A_0_), .B(n2696), .Z(sub_128_aco_B_0_) );
  OR2 C504 ( .A(sub_127_aco_A_10_), .B(sub_127_aco_A_11_), .Z(n2699) );
  OR2 C5051 ( .A(sub_127_aco_A_9_), .B(n2699), .Z(n2700) );
  OR2 C5061 ( .A(sub_127_aco_A_8_), .B(n2700), .Z(n2701) );
  OR2 C5072 ( .A(sub_127_aco_A_7_), .B(n2701), .Z(n2702) );
  OR2 C5081 ( .A(sub_127_aco_A_6_), .B(n2702), .Z(n2703) );
  OR2 C5092 ( .A(sub_127_aco_A_5_), .B(n2703), .Z(n2704) );
  OR2 C5101 ( .A(sub_127_aco_A_4_), .B(n2704), .Z(n2705) );
  OR2 C5112 ( .A(sub_127_aco_A_3_), .B(n2705), .Z(n2706) );
  OR2 C5121 ( .A(sub_127_aco_A_2_), .B(n2706), .Z(n2707) );
  OR2 C5131 ( .A(sub_127_aco_A_1_), .B(n2707), .Z(n2708) );
  OR2 C514 ( .A(sub_127_aco_A_0_), .B(n2708), .Z(sub_127_aco_B_0_) );
  OR2 C5162 ( .A(U3_U1_DATA3_9), .B(U3_U1_DATA3_10), .Z(n2711) );
  OR2 C5172 ( .A(U3_U1_DATA3_8), .B(n2711), .Z(n2712) );
  OR2 C5182 ( .A(U3_U1_DATA3_7), .B(n2712), .Z(n2713) );
  OR2 C5192 ( .A(U3_U1_DATA3_6), .B(n2713), .Z(n2714) );
  OR2 C5202 ( .A(U3_U1_DATA3_5), .B(n2714), .Z(n2715) );
  OR2 C5212 ( .A(U3_U1_DATA3_4), .B(n2715), .Z(n2716) );
  OR2 C5221 ( .A(U3_U1_DATA3_3), .B(n2716), .Z(n2717) );
  OR2 C5231 ( .A(U3_U1_DATA3_2), .B(n2717), .Z(n2718) );
  OR2 C5241 ( .A(U3_U1_DATA3_1), .B(n2718), .Z(n2719) );
  OR2 C5251 ( .A(U3_U1_DATA3_0), .B(n2719), .Z(sub_125_aco_B_0_) );
  OR2 C5271 ( .A(sub_126_aco_A_18_), .B(sub_126_aco_A_19_), .Z(n2722) );
  OR2 C5281 ( .A(sub_126_aco_A_17_), .B(n2722), .Z(n2723) );
  OR2 C5291 ( .A(sub_126_aco_A_16_), .B(n2723), .Z(n2724) );
  OR2 C5302 ( .A(sub_126_aco_A_15_), .B(n2724), .Z(n2725) );
  OR2 C5312 ( .A(sub_126_aco_A_14_), .B(n2725), .Z(n2726) );
  OR2 C5322 ( .A(sub_126_aco_A_13_), .B(n2726), .Z(n2727) );
  OR2 C5332 ( .A(sub_126_aco_A_12_), .B(n2727), .Z(n2728) );
  OR2 C5342 ( .A(sub_126_aco_A_11_), .B(n2728), .Z(n2729) );
  OR2 C5352 ( .A(sub_126_aco_A_10_), .B(n2729), .Z(n2730) );
  OR2 C5362 ( .A(sub_126_aco_A_9_), .B(n2730), .Z(n2731) );
  OR2 C5371 ( .A(sub_126_aco_A_8_), .B(n2731), .Z(n2732) );
  OR2 C5381 ( .A(sub_126_aco_A_7_), .B(n2732), .Z(n2733) );
  OR2 C5392 ( .A(sub_126_aco_A_6_), .B(n2733), .Z(n2734) );
  OR2 C5402 ( .A(sub_126_aco_A_5_), .B(n2734), .Z(n2735) );
  OR2 C5412 ( .A(sub_126_aco_A_4_), .B(n2735), .Z(n2736) );
  OR2 C5421 ( .A(sub_126_aco_A_3_), .B(n2736), .Z(n2737) );
  OR2 C5431 ( .A(sub_126_aco_A_2_), .B(n2737), .Z(n2738) );
  OR2 C5441 ( .A(sub_126_aco_A_1_), .B(n2738), .Z(n2739) );
  OR2 C5451 ( .A(sub_126_aco_A_0_), .B(n2739), .Z(sub_126_aco_B_0_) );
  OR2 C565 ( .A(U76_DATA4_0), .B(n4894), .Z(n2747) );
  OR2 C5811 ( .A(n3273), .B(n4898), .Z(n2749) );
  OR2 C5922 ( .A(U72_DATA2_0), .B(n2593), .Z(n2753) );
  OR2 C5981 ( .A(n2593), .B(n4899), .Z(n2756) );
  OR2 C6031 ( .A(U72_DATA2_0), .B(n4899), .Z(n2757) );
  OR2 C6101 ( .A(n5482), .B(n2587), .Z(n2760) );
  OR2 C6131 ( .A(U76_DATA3_0), .B(U69_DATA4_0), .Z(n2762) );
  OR2 C6421 ( .A(U69_DATA2_0), .B(U71_DATA3_0), .Z(n2770) );
  OR2 C6461 ( .A(U69_DATA2_0), .B(n4903), .Z(n2771) );
  OR2 C655 ( .A(n2774), .B(n2760), .Z(n2775) );
  IV I_1012 ( .A(enable_alternate_refresh), .Z(n2516) );
  OR2 C774 ( .A(n5559), .B(n3273), .Z(n2517) );
  OR2 C814 ( .A(n5481), .B(n2792), .Z(n2587) );
  OR2 C8161 ( .A(n5480), .B(n2791), .Z(n2792) );
  OR2 C8181 ( .A(n5479), .B(n2790), .Z(n2791) );
  OR2 C8201 ( .A(n5478), .B(n2789), .Z(n2790) );
  OR2 C822 ( .A(n5521), .B(n2788), .Z(n2789) );
  OR2 C824 ( .A(n5520), .B(n2787), .Z(n2788) );
  OR2 C8261 ( .A(n5519), .B(n5518), .Z(n2787) );
  AN2 C8421 ( .A(n2793), .B(n5538), .Z(U72_DATA2_0) );
  AN2 C8431 ( .A(n2516), .B(n4900), .Z(n2793) );
  AN2 C8441 ( .A(n2794), .B(n5485), .Z(n2593) );
  AN2 C8451 ( .A(enable_alternate_refresh), .B(n4900), .Z(n2794) );
  AN2 C8511 ( .A(n4900), .B(n5538), .Z(U72_DATA3_0) );
  AN2 C8571 ( .A(n2516), .B(n2517), .Z(U69_DATA2_0) );
  AN2 C858 ( .A(enable_alternate_refresh), .B(n5485), .Z(U71_DATA3_0) );
  AN2 C8681 ( .A(n2795), .B(n5685), .Z(U76_DATA3_0) );
  AN2 C8691 ( .A(n4900), .B(n5572), .Z(n2795) );
  AN2 C8701 ( .A(n5572), .B(n4475), .Z(U69_DATA4_0) );
  AN2 C871 ( .A(n2796), .B(n5685), .Z(U73_DATA5_0) );
  AN2 C872 ( .A(n3273), .B(n5572), .Z(n2796) );
  AN2 C8791 ( .A(n4900), .B(n5582), .Z(U76_DATA4_0) );
  AN2 C8801 ( .A(n3273), .B(n5582), .Z(U73_DATA6_0) );
  IV I_381 ( .A(reset_to_pma_tx), .Z(n2664) );
  AN2 C81 ( .A(n5471), .B(n5470), .Z(n2861) );
  AN2 C91 ( .A(n5469), .B(n5467), .Z(n2862) );
  OR2 C131 ( .A(n5471), .B(U151_DATA3_0), .Z(n2863) );
  OR2 C141 ( .A(U152_DATA3_0), .B(n5467), .Z(n2864) );
  OR2 C191 ( .A(U150_DATA3_0), .B(U151_DATA3_0), .Z(n2867) );
  OR2 C201 ( .A(n5469), .B(n5467), .Z(n2868) );
  OR2 C251 ( .A(n5471), .B(n5470), .Z(n2871) );
  OR2 C261 ( .A(U152_DATA3_0), .B(U153_DATA2_0), .Z(n2872) );
  OR2 C311 ( .A(U150_DATA3_0), .B(n5470), .Z(n2875) );
  OR2 C321 ( .A(U152_DATA3_0), .B(n5467), .Z(n2876) );
  OR2 C372 ( .A(U150_DATA3_0), .B(n5470), .Z(n2879) );
  OR2 C381 ( .A(n5469), .B(U153_DATA2_0), .Z(n2880) );
  OR2 C221 ( .A(U160_DATA2_2), .B(n4921), .Z(n2946) );
  OR2 C222 ( .A(n4918), .B(n2946), .Z(n2947) );
  OR2 C223 ( .A(U160_DATA2_0), .B(n2947), .Z(n2948) );
  OR2 C227 ( .A(n4913), .B(U160_DATA2_3), .Z(n2951) );
  OR2 C228 ( .A(n4918), .B(n2951), .Z(n2952) );
  OR2 C229 ( .A(U160_DATA2_0), .B(n2952), .Z(n2953) );
  OR2 C233 ( .A(U160_DATA2_2), .B(U160_DATA2_3), .Z(n2956) );
  OR2 C234 ( .A(n4918), .B(n2956), .Z(n2957) );
  OR2 C235 ( .A(n4917), .B(n2957), .Z(n2958) );
  OR2 C270 ( .A(U160_DATA2_1), .B(n2946), .Z(n2960) );
  OR2 C2711 ( .A(n4917), .B(n2960), .Z(n2961) );
  OR2 C282 ( .A(U160_DATA2_1), .B(n2951), .Z(n2963) );
  OR2 C283 ( .A(n4917), .B(n2963), .Z(n2964) );
  OR2 C299 ( .A(n4913), .B(n4921), .Z(n2966) );
  OR2 C300 ( .A(U160_DATA2_1), .B(n2966), .Z(n2967) );
  OR2 C301 ( .A(U160_DATA2_0), .B(n2967), .Z(n2968) );
  OR2 C439 ( .A(n2900), .B(U140_CONTROL2), .Z(n2972) );
  OR2 C444 ( .A(n4909), .B(n4915), .Z(n2974) );
  OR2 C4461 ( .A(n4912), .B(U122_CONTROL2), .Z(n2975) );
  OR2 C4501 ( .A(n2892), .B(n4912), .Z(n2977) );
  OR2 C453 ( .A(n2900), .B(U141_CONTROL2), .Z(n2979) );
  OR2 C4661 ( .A(n4916), .B(n4912), .Z(n2985) );
  OR2 C474 ( .A(n4914), .B(n4912), .Z(n2987) );
  OR2 C4761 ( .A(U124_CONTROL2), .B(U122_CONTROL2), .Z(n2988) );
  OR2 C5841 ( .A(n3005), .B(n4912), .Z(n2884) );
  OR2 C5851 ( .A(n3004), .B(n4909), .Z(n3005) );
  OR2 C5861 ( .A(n4911), .B(n4914), .Z(n3004) );
  OR2 C5921 ( .A(n3006), .B(n4909), .Z(n2892) );
  OR2 C5931 ( .A(n4911), .B(n4914), .Z(n3006) );
  OR2 C6001 ( .A(n3008), .B(n4912), .Z(n2900) );
  OR2 C6011 ( .A(n3007), .B(n4916), .Z(n3008) );
  OR2 C6021 ( .A(n4911), .B(n4915), .Z(n3007) );
  OR2 C6141 ( .A(n4911), .B(n4916), .Z(n2915) );
  OR2 C6211 ( .A(n3010), .B(n4909), .Z(n2923) );
  OR2 C6221 ( .A(n3009), .B(n4916), .Z(n3010) );
  OR2 C6231 ( .A(n4911), .B(n4914), .Z(n3009) );
  IV I_281 ( .A(reset_to_pma_tx), .Z(n2937) );
  OR2 C369 ( .A(n4913), .B(U160_DATA2_3), .Z(n3271) );
  OR2 C370 ( .A(n4918), .B(n3271), .Z(n3272) );
  OR2 C371 ( .A(U160_DATA2_0), .B(n3272), .Z(n3273) );
  OR2 C377 ( .A(n5474), .B(tx_mode[1]), .Z(n3279) );
  OR2 C380 ( .A(n5474), .B(tx_mode[1]), .Z(n3281) );
  OR2 C383 ( .A(U149_DATA2_0), .B(n5462), .Z(n3284) );
  OR2 C386 ( .A(n5459), .B(U148_DATA3_0), .Z(n3286) );
  OR2 C389 ( .A(U149_DATA2_0), .B(n5462), .Z(n3288) );
  OR2 C392 ( .A(n5459), .B(U148_DATA3_0), .Z(n3290) );
  OR2 C401 ( .A(n4974), .B(n4949), .Z(n3299) );
  OR2 C402 ( .A(n4997), .B(n3299), .Z(n3300) );
  OR2 C403 ( .A(n5020), .B(n3300), .Z(n3301) );
  OR2 C404 ( .A(n5058), .B(n3301), .Z(n3302) );
  OR2 C405 ( .A(n5081), .B(n3302), .Z(n3303) );
  OR2 C406 ( .A(U162_Z_1), .B(n3303), .Z(n3304) );
  OR2 C407 ( .A(n5093), .B(n3304), .Z(n3305) );
  OR2 C416 ( .A(n5087), .B(n5086), .Z(n3314) );
  OR2 C417 ( .A(n5088), .B(n3314), .Z(n3315) );
  OR2 C418 ( .A(n5089), .B(n3315), .Z(n3316) );
  OR2 C419 ( .A(n5090), .B(n3316), .Z(n3317) );
  OR2 C420 ( .A(n5091), .B(n3317), .Z(n3318) );
  OR2 C421 ( .A(U162_Z_9), .B(n3318), .Z(n3319) );
  OR2 C422 ( .A(n4941), .B(n3319), .Z(n3320) );
  OR2 C431 ( .A(n5078), .B(n5070), .Z(n3329) );
  OR2 C432 ( .A(n5079), .B(n3329), .Z(n3330) );
  OR2 C433 ( .A(n5080), .B(n3330), .Z(n3331) );
  OR2 C434 ( .A(n5082), .B(n3331), .Z(n3332) );
  OR2 C435 ( .A(n5083), .B(n3332), .Z(n3333) );
  OR2 C436 ( .A(U162_Z_17), .B(n3333), .Z(n3334) );
  OR2 C437 ( .A(n5085), .B(n3334), .Z(n3335) );
  OR2 C446 ( .A(n5037), .B(n5028), .Z(n3344) );
  OR2 C447 ( .A(n5038), .B(n3344), .Z(n3345) );
  OR2 C448 ( .A(n5039), .B(n3345), .Z(n3346) );
  OR2 C449 ( .A(n5040), .B(n3346), .Z(n3347) );
  OR2 C450 ( .A(n5041), .B(n3347), .Z(n3348) );
  OR2 C451 ( .A(U162_Z_33), .B(n3348), .Z(n3349) );
  OR2 C452 ( .A(n5043), .B(n3349), .Z(n3350) );
  OR2 C461 ( .A(n5013), .B(n5005), .Z(n3359) );
  OR2 C462 ( .A(n5014), .B(n3359), .Z(n3360) );
  OR2 C463 ( .A(n5015), .B(n3360), .Z(n3361) );
  OR2 C464 ( .A(n5016), .B(n3361), .Z(n3362) );
  OR2 C465 ( .A(n5017), .B(n3362), .Z(n3363) );
  OR2 C466 ( .A(U162_Z_41), .B(n3363), .Z(n3364) );
  OR2 C467 ( .A(n5019), .B(n3364), .Z(n3365) );
  OR2 C476 ( .A(n4992), .B(n4984), .Z(n3374) );
  OR2 C477 ( .A(n4993), .B(n3374), .Z(n3375) );
  OR2 C478 ( .A(n4994), .B(n3375), .Z(n3376) );
  OR2 C479 ( .A(n4995), .B(n3376), .Z(n3377) );
  OR2 C480 ( .A(n4996), .B(n3377), .Z(n3378) );
  OR2 C481 ( .A(U162_Z_49), .B(n3378), .Z(n3379) );
  OR2 C482 ( .A(n4999), .B(n3379), .Z(n3380) );
  OR2 C491 ( .A(n4971), .B(n4963), .Z(n3389) );
  OR2 C492 ( .A(n4972), .B(n3389), .Z(n3390) );
  OR2 C493 ( .A(n4973), .B(n3390), .Z(n3391) );
  OR2 C494 ( .A(n4975), .B(n3391), .Z(n3392) );
  OR2 C495 ( .A(n4976), .B(n3392), .Z(n3393) );
  OR2 C496 ( .A(U162_Z_57), .B(n3393), .Z(n3394) );
  OR2 C497 ( .A(n4978), .B(n3394), .Z(n3395) );
  OR2 C506 ( .A(n5057), .B(n5049), .Z(n3404) );
  OR2 C507 ( .A(n5059), .B(n3404), .Z(n3405) );
  OR2 C508 ( .A(n5060), .B(n3405), .Z(n3406) );
  OR2 C509 ( .A(n5061), .B(n3406), .Z(n3407) );
  OR2 C510 ( .A(n5062), .B(n3407), .Z(n3408) );
  OR2 C511 ( .A(U162_Z_25), .B(n3408), .Z(n3409) );
  OR2 C512 ( .A(n5064), .B(n3409), .Z(n3410) );
  OR2 C515 ( .A(U161_Z_6), .B(U161_Z_7), .Z(n3413) );
  OR2 C516 ( .A(U161_Z_5), .B(n3413), .Z(n3414) );
  OR2 C517 ( .A(U161_Z_4), .B(n3414), .Z(n3415) );
  OR2 C518 ( .A(U161_Z_3), .B(n3415), .Z(n3416) );
  OR2 C519 ( .A(U161_Z_2), .B(n3416), .Z(n3417) );
  OR2 C520 ( .A(U161_Z_1), .B(n3417), .Z(n3418) );
  OR2 C521 ( .A(n5105), .B(n3418), .Z(n3419) );
  OR2 C530 ( .A(n4974), .B(n4949), .Z(n3422) );
  OR2 C531 ( .A(n4997), .B(n3422), .Z(n3423) );
  OR2 C532 ( .A(n5020), .B(n3423), .Z(n3424) );
  OR2 C533 ( .A(n5058), .B(n3424), .Z(n3425) );
  OR2 C534 ( .A(U162_Z_2), .B(n3425), .Z(n3426) );
  OR2 C535 ( .A(n5092), .B(n3426), .Z(n3427) );
  OR2 C536 ( .A(n5093), .B(n3427), .Z(n3428) );
  OR2 C539 ( .A(U161_Z_6), .B(U161_Z_7), .Z(n3431) );
  OR2 C540 ( .A(U161_Z_5), .B(n3431), .Z(n3432) );
  OR2 C541 ( .A(n5100), .B(n3432), .Z(n3433) );
  OR2 C550 ( .A(n5037), .B(n5028), .Z(n3436) );
  OR2 C551 ( .A(n5038), .B(n3436), .Z(n3437) );
  OR2 C552 ( .A(n5039), .B(n3437), .Z(n3438) );
  OR2 C553 ( .A(n5040), .B(n3438), .Z(n3439) );
  OR2 C554 ( .A(U162_Z_34), .B(n3439), .Z(n3440) );
  OR2 C555 ( .A(n5042), .B(n3440), .Z(n3441) );
  OR2 C556 ( .A(n5043), .B(n3441), .Z(n3442) );
  OR2 C558 ( .A(n3218), .B(n3217), .Z(n3444) );
  OR2 C559 ( .A(n3219), .B(n3444), .Z(n3445) );
  OR2 C560 ( .A(n3220), .B(n3445), .Z(n3446) );
  OR2 C561 ( .A(n3221), .B(n3446), .Z(n3447) );
  OR2 C562 ( .A(n3222), .B(n3447), .Z(n3448) );
  OR2 C563 ( .A(n3223), .B(n3448), .Z(n3449) );
  OR2 C564 ( .A(n3224), .B(n3449), .Z(n3450) );
  OR2 C570 ( .A(n4990), .B(n4969), .Z(n3456) );
  OR2 C571 ( .A(n5011), .B(n3456), .Z(n3457) );
  OR2 C572 ( .A(n5034), .B(n3457), .Z(n3458) );
  OR2 C573 ( .A(n3221), .B(n3458), .Z(n3459) );
  OR2 C574 ( .A(n3222), .B(n3459), .Z(n3460) );
  OR2 C575 ( .A(n3223), .B(n3460), .Z(n3461) );
  OR2 C576 ( .A(n3224), .B(n3461), .Z(n3462) );
  OR2 C582 ( .A(n3218), .B(n3217), .Z(n3468) );
  OR2 C583 ( .A(n3219), .B(n3468), .Z(n3469) );
  OR2 C584 ( .A(n3220), .B(n3469), .Z(n3470) );
  OR2 C585 ( .A(n5055), .B(n3470), .Z(n3471) );
  OR2 C586 ( .A(n5076), .B(n3471), .Z(n3472) );
  OR2 C587 ( .A(n4929), .B(n3472), .Z(n3473) );
  OR2 C588 ( .A(n4955), .B(n3473), .Z(n3474) );
  IV I_96 ( .A(tx_fifo_pop_pre), .Z(n3476) );
  OR2 C592 ( .A(U161_Z_2), .B(U161_Z_3), .Z(n3477) );
  OR2 C593 ( .A(U161_Z_1), .B(n3477), .Z(n3478) );
  OR2 C594 ( .A(n5105), .B(n3478), .Z(n3479) );
  OR2 C600 ( .A(U162_Z_6), .B(n4949), .Z(n3481) );
  OR2 C601 ( .A(U162_Z_5), .B(n3481), .Z(n3482) );
  OR2 C602 ( .A(n5020), .B(n3482), .Z(n3483) );
  OR2 C603 ( .A(n5058), .B(n3483), .Z(n3484) );
  OR2 C604 ( .A(n5081), .B(n3484), .Z(n3485) );
  OR2 C605 ( .A(U162_Z_1), .B(n3485), .Z(n3486) );
  OR2 C606 ( .A(U162_Z_0), .B(n3486), .Z(n3487) );
  OR2 C612 ( .A(n4974), .B(U162_Z_7), .Z(n3489) );
  OR2 C613 ( .A(U162_Z_5), .B(n3489), .Z(n3490) );
  OR2 C614 ( .A(n5020), .B(n3490), .Z(n3491) );
  OR2 C615 ( .A(n5058), .B(n3491), .Z(n3492) );
  OR2 C616 ( .A(n5081), .B(n3492), .Z(n3493) );
  OR2 C617 ( .A(U162_Z_1), .B(n3493), .Z(n3494) );
  OR2 C618 ( .A(U162_Z_0), .B(n3494), .Z(n3495) );
  OR2 C621 ( .A(U161_Z_6), .B(U161_Z_7), .Z(n3497) );
  OR2 C622 ( .A(U161_Z_5), .B(n3497), .Z(n3498) );
  OR2 C623 ( .A(n5100), .B(n3498), .Z(n3499) );
  OR2 C629 ( .A(U162_Z_38), .B(n5028), .Z(n3501) );
  OR2 C630 ( .A(U162_Z_37), .B(n3501), .Z(n3502) );
  OR2 C631 ( .A(n5039), .B(n3502), .Z(n3503) );
  OR2 C632 ( .A(n5040), .B(n3503), .Z(n3504) );
  OR2 C633 ( .A(n5041), .B(n3504), .Z(n3505) );
  OR2 C634 ( .A(U162_Z_33), .B(n3505), .Z(n3506) );
  OR2 C635 ( .A(U162_Z_32), .B(n3506), .Z(n3507) );
  OR2 C641 ( .A(n5037), .B(U162_Z_39), .Z(n3509) );
  OR2 C642 ( .A(U162_Z_37), .B(n3509), .Z(n3510) );
  OR2 C643 ( .A(n5039), .B(n3510), .Z(n3511) );
  OR2 C644 ( .A(n5040), .B(n3511), .Z(n3512) );
  OR2 C645 ( .A(n5041), .B(n3512), .Z(n3513) );
  OR2 C646 ( .A(U162_Z_33), .B(n3513), .Z(n3514) );
  OR2 C647 ( .A(U162_Z_32), .B(n3514), .Z(n3515) );
  OR2 C651 ( .A(n5455), .B(n[3181]), .Z(n3519) );
  OR2 C652 ( .A(n5454), .B(n3519), .Z(n3520) );
  OR2 C653 ( .A(n[3184]), .B(n3520), .Z(n3521) );
  OR2 C657 ( .A(U162_Z_6), .B(U162_Z_7), .Z(n3523) );
  OR2 C658 ( .A(U162_Z_5), .B(n3523), .Z(n3524) );
  OR2 C659 ( .A(U162_Z_4), .B(n3524), .Z(n3525) );
  OR2 C660 ( .A(U162_Z_3), .B(n3525), .Z(n3526) );
  OR2 C661 ( .A(n5081), .B(n3526), .Z(n3527) );
  OR2 C662 ( .A(n5092), .B(n3527), .Z(n3528) );
  OR2 C663 ( .A(U162_Z_0), .B(n3528), .Z(n3529) );
  OR2 C667 ( .A(U162_Z_14), .B(U162_Z_15), .Z(n3532) );
  OR2 C668 ( .A(U162_Z_13), .B(n3532), .Z(n3533) );
  OR2 C669 ( .A(U162_Z_12), .B(n3533), .Z(n3534) );
  OR2 C670 ( .A(U162_Z_11), .B(n3534), .Z(n3535) );
  OR2 C671 ( .A(n5091), .B(n3535), .Z(n3536) );
  OR2 C672 ( .A(n4934), .B(n3536), .Z(n3537) );
  OR2 C673 ( .A(U162_Z_8), .B(n3537), .Z(n3538) );
  OR2 C677 ( .A(U162_Z_22), .B(U162_Z_23), .Z(n3541) );
  OR2 C678 ( .A(U162_Z_21), .B(n3541), .Z(n3542) );
  OR2 C679 ( .A(U162_Z_20), .B(n3542), .Z(n3543) );
  OR2 C680 ( .A(U162_Z_19), .B(n3543), .Z(n3544) );
  OR2 C681 ( .A(n5083), .B(n3544), .Z(n3545) );
  OR2 C682 ( .A(n5084), .B(n3545), .Z(n3546) );
  OR2 C683 ( .A(U162_Z_16), .B(n3546), .Z(n3547) );
  OR2 C687 ( .A(U162_Z_30), .B(U162_Z_31), .Z(n3550) );
  OR2 C688 ( .A(U162_Z_29), .B(n3550), .Z(n3551) );
  OR2 C689 ( .A(U162_Z_28), .B(n3551), .Z(n3552) );
  OR2 C690 ( .A(U162_Z_27), .B(n3552), .Z(n3553) );
  OR2 C691 ( .A(n5062), .B(n3553), .Z(n3554) );
  OR2 C692 ( .A(n5063), .B(n3554), .Z(n3555) );
  OR2 C693 ( .A(U162_Z_24), .B(n3555), .Z(n3556) );
  OR2 C697 ( .A(U162_Z_38), .B(U162_Z_39), .Z(n3558) );
  OR2 C698 ( .A(U162_Z_37), .B(n3558), .Z(n3559) );
  OR2 C699 ( .A(U162_Z_36), .B(n3559), .Z(n3560) );
  OR2 C700 ( .A(U162_Z_35), .B(n3560), .Z(n3561) );
  OR2 C701 ( .A(n5041), .B(n3561), .Z(n3562) );
  OR2 C702 ( .A(n5042), .B(n3562), .Z(n3563) );
  OR2 C703 ( .A(U162_Z_32), .B(n3563), .Z(n3564) );
  OR2 C707 ( .A(U162_Z_46), .B(U162_Z_47), .Z(n3567) );
  OR2 C708 ( .A(U162_Z_45), .B(n3567), .Z(n3568) );
  OR2 C709 ( .A(U162_Z_44), .B(n3568), .Z(n3569) );
  OR2 C710 ( .A(U162_Z_43), .B(n3569), .Z(n3570) );
  OR2 C711 ( .A(n5017), .B(n3570), .Z(n3571) );
  OR2 C712 ( .A(n5018), .B(n3571), .Z(n3572) );
  OR2 C713 ( .A(U162_Z_40), .B(n3572), .Z(n3573) );
  OR2 C717 ( .A(U162_Z_54), .B(U162_Z_55), .Z(n3576) );
  OR2 C718 ( .A(U162_Z_53), .B(n3576), .Z(n3577) );
  OR2 C719 ( .A(U162_Z_52), .B(n3577), .Z(n3578) );
  OR2 C720 ( .A(U162_Z_51), .B(n3578), .Z(n3579) );
  OR2 C721 ( .A(n4996), .B(n3579), .Z(n3580) );
  OR2 C722 ( .A(n4998), .B(n3580), .Z(n3581) );
  OR2 C723 ( .A(U162_Z_48), .B(n3581), .Z(n3582) );
  OR2 C727 ( .A(U162_Z_62), .B(U162_Z_63), .Z(n3585) );
  OR2 C728 ( .A(U162_Z_61), .B(n3585), .Z(n3586) );
  OR2 C729 ( .A(U162_Z_60), .B(n3586), .Z(n3587) );
  OR2 C730 ( .A(U162_Z_59), .B(n3587), .Z(n3588) );
  OR2 C731 ( .A(n4976), .B(n3588), .Z(n3589) );
  OR2 C732 ( .A(n4977), .B(n3589), .Z(n3590) );
  OR2 C733 ( .A(U162_Z_56), .B(n3590), .Z(n3591) );
  OR2 C738 ( .A(U162_Z_38), .B(U162_Z_39), .Z(n3593) );
  OR2 C739 ( .A(U162_Z_37), .B(n3593), .Z(n3594) );
  OR2 C740 ( .A(U162_Z_36), .B(n3594), .Z(n3595) );
  OR2 C741 ( .A(U162_Z_35), .B(n3595), .Z(n3596) );
  OR2 C742 ( .A(n5041), .B(n3596), .Z(n3597) );
  OR2 C743 ( .A(n5042), .B(n3597), .Z(n3598) );
  OR2 C744 ( .A(n5043), .B(n3598), .Z(n3599) );
  OR2 C751 ( .A(n5037), .B(U162_Z_39), .Z(n3601) );
  OR2 C752 ( .A(n5038), .B(n3601), .Z(n3602) );
  OR2 C753 ( .A(n5039), .B(n3602), .Z(n3603) );
  OR2 C754 ( .A(n5040), .B(n3603), .Z(n3604) );
  OR2 C755 ( .A(n5041), .B(n3604), .Z(n3605) );
  OR2 C756 ( .A(U162_Z_33), .B(n3605), .Z(n3606) );
  OR2 C757 ( .A(U162_Z_32), .B(n3606), .Z(n3607) );
  OR2 C762 ( .A(U162_Z_38), .B(U162_Z_39), .Z(n3609) );
  OR2 C763 ( .A(U162_Z_37), .B(n3609), .Z(n3610) );
  OR2 C764 ( .A(n5039), .B(n3610), .Z(n3611) );
  OR2 C765 ( .A(n5040), .B(n3611), .Z(n3612) );
  OR2 C766 ( .A(n5041), .B(n3612), .Z(n3613) );
  OR2 C767 ( .A(U162_Z_33), .B(n3613), .Z(n3614) );
  OR2 C768 ( .A(U162_Z_32), .B(n3614), .Z(n3615) );
  OR2 C775 ( .A(U162_Z_38), .B(n5028), .Z(n3617) );
  OR2 C776 ( .A(n5038), .B(n3617), .Z(n3618) );
  OR2 C777 ( .A(n5039), .B(n3618), .Z(n3619) );
  OR2 C778 ( .A(n5040), .B(n3619), .Z(n3620) );
  OR2 C779 ( .A(n5041), .B(n3620), .Z(n3621) );
  OR2 C780 ( .A(U162_Z_33), .B(n3621), .Z(n3622) );
  OR2 C781 ( .A(U162_Z_32), .B(n3622), .Z(n3623) );
  OR2 C787 ( .A(U162_Z_38), .B(U162_Z_39), .Z(n3625) );
  OR2 C788 ( .A(n5038), .B(n3625), .Z(n3626) );
  OR2 C789 ( .A(n5039), .B(n3626), .Z(n3627) );
  OR2 C790 ( .A(n5040), .B(n3627), .Z(n3628) );
  OR2 C791 ( .A(n5041), .B(n3628), .Z(n3629) );
  OR2 C792 ( .A(U162_Z_33), .B(n3629), .Z(n3630) );
  OR2 C793 ( .A(U162_Z_32), .B(n3630), .Z(n3631) );
  OR2 C800 ( .A(n5037), .B(n5028), .Z(n3633) );
  OR2 C801 ( .A(U162_Z_37), .B(n3633), .Z(n3634) );
  OR2 C802 ( .A(n5039), .B(n3634), .Z(n3635) );
  OR2 C803 ( .A(n5040), .B(n3635), .Z(n3636) );
  OR2 C804 ( .A(n5041), .B(n3636), .Z(n3637) );
  OR2 C805 ( .A(U162_Z_33), .B(n3637), .Z(n3638) );
  OR2 C806 ( .A(U162_Z_32), .B(n3638), .Z(n3639) );
  OR2 C815 ( .A(n5037), .B(n5028), .Z(n3641) );
  OR2 C816 ( .A(n5038), .B(n3641), .Z(n3642) );
  OR2 C817 ( .A(n5039), .B(n3642), .Z(n3643) );
  OR2 C818 ( .A(U162_Z_35), .B(n3643), .Z(n3644) );
  OR2 C819 ( .A(n5041), .B(n3644), .Z(n3645) );
  OR2 C820 ( .A(n5042), .B(n3645), .Z(n3646) );
  OR2 C821 ( .A(n5043), .B(n3646), .Z(n3647) );
  OR2 C825 ( .A(U162_Z_38), .B(U162_Z_39), .Z(n3649) );
  OR2 C826 ( .A(U162_Z_37), .B(n3649), .Z(n3650) );
  OR2 C827 ( .A(U162_Z_36), .B(n3650), .Z(n3651) );
  OR2 C828 ( .A(U162_Z_35), .B(n3651), .Z(n3652) );
  OR2 C829 ( .A(n5041), .B(n3652), .Z(n3653) );
  OR2 C830 ( .A(n5042), .B(n3653), .Z(n3654) );
  OR2 C831 ( .A(U162_Z_32), .B(n3654), .Z(n3655) );
  OR2 C840 ( .A(n5037), .B(n5028), .Z(n3657) );
  OR2 C841 ( .A(n5038), .B(n3657), .Z(n3658) );
  OR2 C842 ( .A(n5039), .B(n3658), .Z(n3659) );
  OR2 C843 ( .A(n5040), .B(n3659), .Z(n3660) );
  OR2 C844 ( .A(n5041), .B(n3660), .Z(n3661) );
  OR2 C845 ( .A(n5042), .B(n3661), .Z(n3662) );
  OR2 C846 ( .A(U162_Z_32), .B(n3662), .Z(n3663) );
  OR2 C851 ( .A(U162_Z_46), .B(U162_Z_47), .Z(n3665) );
  OR2 C852 ( .A(U162_Z_45), .B(n3665), .Z(n3666) );
  OR2 C853 ( .A(U162_Z_44), .B(n3666), .Z(n3667) );
  OR2 C854 ( .A(U162_Z_43), .B(n3667), .Z(n3668) );
  OR2 C855 ( .A(n5017), .B(n3668), .Z(n3669) );
  OR2 C856 ( .A(n5018), .B(n3669), .Z(n3670) );
  OR2 C857 ( .A(n5019), .B(n3670), .Z(n3671) );
  OR2 C864 ( .A(n5013), .B(U162_Z_47), .Z(n3673) );
  OR2 C865 ( .A(n5014), .B(n3673), .Z(n3674) );
  OR2 C866 ( .A(n5015), .B(n3674), .Z(n3675) );
  OR2 C867 ( .A(n5016), .B(n3675), .Z(n3676) );
  OR2 C868 ( .A(n5017), .B(n3676), .Z(n3677) );
  OR2 C869 ( .A(U162_Z_41), .B(n3677), .Z(n3678) );
  OR2 C870 ( .A(U162_Z_40), .B(n3678), .Z(n3679) );
  OR2 C875 ( .A(U162_Z_46), .B(U162_Z_47), .Z(n3681) );
  OR2 C876 ( .A(U162_Z_45), .B(n3681), .Z(n3682) );
  OR2 C877 ( .A(n5015), .B(n3682), .Z(n3683) );
  OR2 C878 ( .A(n5016), .B(n3683), .Z(n3684) );
  OR2 C879 ( .A(n5017), .B(n3684), .Z(n3685) );
  OR2 C880 ( .A(U162_Z_41), .B(n3685), .Z(n3686) );
  OR2 C881 ( .A(U162_Z_40), .B(n3686), .Z(n3687) );
  OR2 C888 ( .A(U162_Z_46), .B(n5005), .Z(n3689) );
  OR2 C889 ( .A(n5014), .B(n3689), .Z(n3690) );
  OR2 C890 ( .A(n5015), .B(n3690), .Z(n3691) );
  OR2 C891 ( .A(n5016), .B(n3691), .Z(n3692) );
  OR2 C892 ( .A(n5017), .B(n3692), .Z(n3693) );
  OR2 C893 ( .A(U162_Z_41), .B(n3693), .Z(n3694) );
  OR2 C894 ( .A(U162_Z_40), .B(n3694), .Z(n3695) );
  OR2 C900 ( .A(U162_Z_46), .B(U162_Z_47), .Z(n3697) );
  OR2 C901 ( .A(n5014), .B(n3697), .Z(n3698) );
  OR2 C902 ( .A(n5015), .B(n3698), .Z(n3699) );
  OR2 C903 ( .A(n5016), .B(n3699), .Z(n3700) );
  OR2 C904 ( .A(n5017), .B(n3700), .Z(n3701) );
  OR2 C905 ( .A(U162_Z_41), .B(n3701), .Z(n3702) );
  OR2 C906 ( .A(U162_Z_40), .B(n3702), .Z(n3703) );
  OR2 C913 ( .A(n5013), .B(n5005), .Z(n3705) );
  OR2 C914 ( .A(U162_Z_45), .B(n3705), .Z(n3706) );
  OR2 C915 ( .A(n5015), .B(n3706), .Z(n3707) );
  OR2 C916 ( .A(n5016), .B(n3707), .Z(n3708) );
  OR2 C917 ( .A(n5017), .B(n3708), .Z(n3709) );
  OR2 C918 ( .A(U162_Z_41), .B(n3709), .Z(n3710) );
  OR2 C919 ( .A(U162_Z_40), .B(n3710), .Z(n3711) );
  OR2 C928 ( .A(n5013), .B(n5005), .Z(n3713) );
  OR2 C929 ( .A(n5014), .B(n3713), .Z(n3714) );
  OR2 C930 ( .A(n5015), .B(n3714), .Z(n3715) );
  OR2 C931 ( .A(U162_Z_43), .B(n3715), .Z(n3716) );
  OR2 C932 ( .A(n5017), .B(n3716), .Z(n3717) );
  OR2 C933 ( .A(n5018), .B(n3717), .Z(n3718) );
  OR2 C934 ( .A(n5019), .B(n3718), .Z(n3719) );
  OR2 C938 ( .A(U162_Z_46), .B(U162_Z_47), .Z(n3721) );
  OR2 C939 ( .A(U162_Z_45), .B(n3721), .Z(n3722) );
  OR2 C940 ( .A(U162_Z_44), .B(n3722), .Z(n3723) );
  OR2 C941 ( .A(U162_Z_43), .B(n3723), .Z(n3724) );
  OR2 C942 ( .A(n5017), .B(n3724), .Z(n3725) );
  OR2 C943 ( .A(n5018), .B(n3725), .Z(n3726) );
  OR2 C944 ( .A(U162_Z_40), .B(n3726), .Z(n3727) );
  OR2 C953 ( .A(n5013), .B(n5005), .Z(n3729) );
  OR2 C954 ( .A(n5014), .B(n3729), .Z(n3730) );
  OR2 C955 ( .A(n5015), .B(n3730), .Z(n3731) );
  OR2 C956 ( .A(n5016), .B(n3731), .Z(n3732) );
  OR2 C957 ( .A(n5017), .B(n3732), .Z(n3733) );
  OR2 C958 ( .A(n5018), .B(n3733), .Z(n3734) );
  OR2 C959 ( .A(U162_Z_40), .B(n3734), .Z(n3735) );
  OR2 C964 ( .A(U162_Z_54), .B(U162_Z_55), .Z(n3737) );
  OR2 C965 ( .A(U162_Z_53), .B(n3737), .Z(n3738) );
  OR2 C966 ( .A(U162_Z_52), .B(n3738), .Z(n3739) );
  OR2 C967 ( .A(U162_Z_51), .B(n3739), .Z(n3740) );
  OR2 C968 ( .A(n4996), .B(n3740), .Z(n3741) );
  OR2 C969 ( .A(n4998), .B(n3741), .Z(n3742) );
  OR2 C970 ( .A(n4999), .B(n3742), .Z(n3743) );
  OR2 C977 ( .A(n4992), .B(U162_Z_55), .Z(n3745) );
  OR2 C978 ( .A(n4993), .B(n3745), .Z(n3746) );
  OR2 C979 ( .A(n4994), .B(n3746), .Z(n3747) );
  OR2 C980 ( .A(n4995), .B(n3747), .Z(n3748) );
  OR2 C981 ( .A(n4996), .B(n3748), .Z(n3749) );
  OR2 C982 ( .A(U162_Z_49), .B(n3749), .Z(n3750) );
  OR2 C983 ( .A(U162_Z_48), .B(n3750), .Z(n3751) );
  OR2 C988 ( .A(U162_Z_54), .B(U162_Z_55), .Z(n3753) );
  OR2 C989 ( .A(U162_Z_53), .B(n3753), .Z(n3754) );
  OR2 C990 ( .A(n4994), .B(n3754), .Z(n3755) );
  OR2 C991 ( .A(n4995), .B(n3755), .Z(n3756) );
  OR2 C992 ( .A(n4996), .B(n3756), .Z(n3757) );
  OR2 C993 ( .A(U162_Z_49), .B(n3757), .Z(n3758) );
  OR2 C994 ( .A(U162_Z_48), .B(n3758), .Z(n3759) );
  OR2 C1001 ( .A(U162_Z_54), .B(n4984), .Z(n3761) );
  OR2 C1002 ( .A(n4993), .B(n3761), .Z(n3762) );
  OR2 C1003 ( .A(n4994), .B(n3762), .Z(n3763) );
  OR2 C1004 ( .A(n4995), .B(n3763), .Z(n3764) );
  OR2 C1005 ( .A(n4996), .B(n3764), .Z(n3765) );
  OR2 C1006 ( .A(U162_Z_49), .B(n3765), .Z(n3766) );
  OR2 C1007 ( .A(U162_Z_48), .B(n3766), .Z(n3767) );
  OR2 C1013 ( .A(U162_Z_54), .B(U162_Z_55), .Z(n3769) );
  OR2 C1014 ( .A(n4993), .B(n3769), .Z(n3770) );
  OR2 C1015 ( .A(n4994), .B(n3770), .Z(n3771) );
  OR2 C1016 ( .A(n4995), .B(n3771), .Z(n3772) );
  OR2 C1017 ( .A(n4996), .B(n3772), .Z(n3773) );
  OR2 C1018 ( .A(U162_Z_49), .B(n3773), .Z(n3774) );
  OR2 C1019 ( .A(U162_Z_48), .B(n3774), .Z(n3775) );
  OR2 C1026 ( .A(n4992), .B(n4984), .Z(n3777) );
  OR2 C1027 ( .A(U162_Z_53), .B(n3777), .Z(n3778) );
  OR2 C1028 ( .A(n4994), .B(n3778), .Z(n3779) );
  OR2 C1029 ( .A(n4995), .B(n3779), .Z(n3780) );
  OR2 C1030 ( .A(n4996), .B(n3780), .Z(n3781) );
  OR2 C1031 ( .A(U162_Z_49), .B(n3781), .Z(n3782) );
  OR2 C1032 ( .A(U162_Z_48), .B(n3782), .Z(n3783) );
  OR2 C1041 ( .A(n4992), .B(n4984), .Z(n3785) );
  OR2 C1042 ( .A(n4993), .B(n3785), .Z(n3786) );
  OR2 C1043 ( .A(n4994), .B(n3786), .Z(n3787) );
  OR2 C1044 ( .A(U162_Z_51), .B(n3787), .Z(n3788) );
  OR2 C1045 ( .A(n4996), .B(n3788), .Z(n3789) );
  OR2 C1046 ( .A(n4998), .B(n3789), .Z(n3790) );
  OR2 C1047 ( .A(n4999), .B(n3790), .Z(n3791) );
  OR2 C1051 ( .A(U162_Z_54), .B(U162_Z_55), .Z(n3793) );
  OR2 C1052 ( .A(U162_Z_53), .B(n3793), .Z(n3794) );
  OR2 C1053 ( .A(U162_Z_52), .B(n3794), .Z(n3795) );
  OR2 C1054 ( .A(U162_Z_51), .B(n3795), .Z(n3796) );
  OR2 C1055 ( .A(n4996), .B(n3796), .Z(n3797) );
  OR2 C1056 ( .A(n4998), .B(n3797), .Z(n3798) );
  OR2 C1057 ( .A(U162_Z_48), .B(n3798), .Z(n3799) );
  OR2 C1066 ( .A(n4992), .B(n4984), .Z(n3801) );
  OR2 C1067 ( .A(n4993), .B(n3801), .Z(n3802) );
  OR2 C1068 ( .A(n4994), .B(n3802), .Z(n3803) );
  OR2 C1069 ( .A(n4995), .B(n3803), .Z(n3804) );
  OR2 C1070 ( .A(n4996), .B(n3804), .Z(n3805) );
  OR2 C1071 ( .A(n4998), .B(n3805), .Z(n3806) );
  OR2 C1072 ( .A(U162_Z_48), .B(n3806), .Z(n3807) );
  OR2 C1077 ( .A(U162_Z_62), .B(U162_Z_63), .Z(n3809) );
  OR2 C1078 ( .A(U162_Z_61), .B(n3809), .Z(n3810) );
  OR2 C1079 ( .A(U162_Z_60), .B(n3810), .Z(n3811) );
  OR2 C1080 ( .A(U162_Z_59), .B(n3811), .Z(n3812) );
  OR2 C1081 ( .A(n4976), .B(n3812), .Z(n3813) );
  OR2 C1082 ( .A(n4977), .B(n3813), .Z(n3814) );
  OR2 C1083 ( .A(n4978), .B(n3814), .Z(n3815) );
  OR2 C1090 ( .A(n4971), .B(U162_Z_63), .Z(n3817) );
  OR2 C1091 ( .A(n4972), .B(n3817), .Z(n3818) );
  OR2 C1092 ( .A(n4973), .B(n3818), .Z(n3819) );
  OR2 C1093 ( .A(n4975), .B(n3819), .Z(n3820) );
  OR2 C1094 ( .A(n4976), .B(n3820), .Z(n3821) );
  OR2 C1095 ( .A(U162_Z_57), .B(n3821), .Z(n3822) );
  OR2 C1096 ( .A(U162_Z_56), .B(n3822), .Z(n3823) );
  OR2 C1101 ( .A(U162_Z_62), .B(U162_Z_63), .Z(n3825) );
  OR2 C1102 ( .A(U162_Z_61), .B(n3825), .Z(n3826) );
  OR2 C1103 ( .A(n4973), .B(n3826), .Z(n3827) );
  OR2 C1104 ( .A(n4975), .B(n3827), .Z(n3828) );
  OR2 C1105 ( .A(n4976), .B(n3828), .Z(n3829) );
  OR2 C1106 ( .A(U162_Z_57), .B(n3829), .Z(n3830) );
  OR2 C1107 ( .A(U162_Z_56), .B(n3830), .Z(n3831) );
  OR2 C1114 ( .A(U162_Z_62), .B(n4963), .Z(n3833) );
  OR2 C1115 ( .A(n4972), .B(n3833), .Z(n3834) );
  OR2 C1116 ( .A(n4973), .B(n3834), .Z(n3835) );
  OR2 C1117 ( .A(n4975), .B(n3835), .Z(n3836) );
  OR2 C1118 ( .A(n4976), .B(n3836), .Z(n3837) );
  OR2 C1119 ( .A(U162_Z_57), .B(n3837), .Z(n3838) );
  OR2 C1120 ( .A(U162_Z_56), .B(n3838), .Z(n3839) );
  OR2 C1126 ( .A(U162_Z_62), .B(U162_Z_63), .Z(n3841) );
  OR2 C1127 ( .A(n4972), .B(n3841), .Z(n3842) );
  OR2 C1128 ( .A(n4973), .B(n3842), .Z(n3843) );
  OR2 C1129 ( .A(n4975), .B(n3843), .Z(n3844) );
  OR2 C1130 ( .A(n4976), .B(n3844), .Z(n3845) );
  OR2 C1131 ( .A(U162_Z_57), .B(n3845), .Z(n3846) );
  OR2 C1132 ( .A(U162_Z_56), .B(n3846), .Z(n3847) );
  OR2 C1139 ( .A(n4971), .B(n4963), .Z(n3849) );
  OR2 C1140 ( .A(U162_Z_61), .B(n3849), .Z(n3850) );
  OR2 C1141 ( .A(n4973), .B(n3850), .Z(n3851) );
  OR2 C1142 ( .A(n4975), .B(n3851), .Z(n3852) );
  OR2 C1143 ( .A(n4976), .B(n3852), .Z(n3853) );
  OR2 C1144 ( .A(U162_Z_57), .B(n3853), .Z(n3854) );
  OR2 C1145 ( .A(U162_Z_56), .B(n3854), .Z(n3855) );
  OR2 C1154 ( .A(n4971), .B(n4963), .Z(n3857) );
  OR2 C1155 ( .A(n4972), .B(n3857), .Z(n3858) );
  OR2 C1156 ( .A(n4973), .B(n3858), .Z(n3859) );
  OR2 C1157 ( .A(U162_Z_59), .B(n3859), .Z(n3860) );
  OR2 C1158 ( .A(n4976), .B(n3860), .Z(n3861) );
  OR2 C1159 ( .A(n4977), .B(n3861), .Z(n3862) );
  OR2 C1160 ( .A(n4978), .B(n3862), .Z(n3863) );
  OR2 C1164 ( .A(U162_Z_62), .B(U162_Z_63), .Z(n3865) );
  OR2 C1165 ( .A(U162_Z_61), .B(n3865), .Z(n3866) );
  OR2 C1166 ( .A(U162_Z_60), .B(n3866), .Z(n3867) );
  OR2 C1167 ( .A(U162_Z_59), .B(n3867), .Z(n3868) );
  OR2 C1168 ( .A(n4976), .B(n3868), .Z(n3869) );
  OR2 C1169 ( .A(n4977), .B(n3869), .Z(n3870) );
  OR2 C1170 ( .A(U162_Z_56), .B(n3870), .Z(n3871) );
  OR2 C1179 ( .A(n4971), .B(n4963), .Z(n3873) );
  OR2 C1180 ( .A(n4972), .B(n3873), .Z(n3874) );
  OR2 C1181 ( .A(n4973), .B(n3874), .Z(n3875) );
  OR2 C1182 ( .A(n4975), .B(n3875), .Z(n3876) );
  OR2 C1183 ( .A(n4976), .B(n3876), .Z(n3877) );
  OR2 C1184 ( .A(n4977), .B(n3877), .Z(n3878) );
  OR2 C1185 ( .A(U162_Z_56), .B(n3878), .Z(n3879) );
  OR2 C1190 ( .A(U162_Z_6), .B(U162_Z_7), .Z(n3881) );
  OR2 C1191 ( .A(U162_Z_5), .B(n3881), .Z(n3882) );
  OR2 C1192 ( .A(U162_Z_4), .B(n3882), .Z(n3883) );
  OR2 C1193 ( .A(U162_Z_3), .B(n3883), .Z(n3884) );
  OR2 C1194 ( .A(n5081), .B(n3884), .Z(n3885) );
  OR2 C1195 ( .A(n5092), .B(n3885), .Z(n3886) );
  OR2 C1196 ( .A(n5093), .B(n3886), .Z(n3887) );
  OR2 C1203 ( .A(n4974), .B(U162_Z_7), .Z(n3889) );
  OR2 C1204 ( .A(n4997), .B(n3889), .Z(n3890) );
  OR2 C1205 ( .A(n5020), .B(n3890), .Z(n3891) );
  OR2 C1206 ( .A(n5058), .B(n3891), .Z(n3892) );
  OR2 C1207 ( .A(n5081), .B(n3892), .Z(n3893) );
  OR2 C1208 ( .A(U162_Z_1), .B(n3893), .Z(n3894) );
  OR2 C1209 ( .A(U162_Z_0), .B(n3894), .Z(n3895) );
  OR2 C1214 ( .A(U162_Z_6), .B(U162_Z_7), .Z(n3897) );
  OR2 C1215 ( .A(U162_Z_5), .B(n3897), .Z(n3898) );
  OR2 C1216 ( .A(n5020), .B(n3898), .Z(n3899) );
  OR2 C1217 ( .A(n5058), .B(n3899), .Z(n3900) );
  OR2 C1218 ( .A(n5081), .B(n3900), .Z(n3901) );
  OR2 C1219 ( .A(U162_Z_1), .B(n3901), .Z(n3902) );
  OR2 C1220 ( .A(U162_Z_0), .B(n3902), .Z(n3903) );
  OR2 C1227 ( .A(U162_Z_6), .B(n4949), .Z(n3905) );
  OR2 C1228 ( .A(n4997), .B(n3905), .Z(n3906) );
  OR2 C1229 ( .A(n5020), .B(n3906), .Z(n3907) );
  OR2 C1230 ( .A(n5058), .B(n3907), .Z(n3908) );
  OR2 C1231 ( .A(n5081), .B(n3908), .Z(n3909) );
  OR2 C1232 ( .A(U162_Z_1), .B(n3909), .Z(n3910) );
  OR2 C1233 ( .A(U162_Z_0), .B(n3910), .Z(n3911) );
  OR2 C1239 ( .A(U162_Z_6), .B(U162_Z_7), .Z(n3913) );
  OR2 C1240 ( .A(n4997), .B(n3913), .Z(n3914) );
  OR2 C1241 ( .A(n5020), .B(n3914), .Z(n3915) );
  OR2 C1242 ( .A(n5058), .B(n3915), .Z(n3916) );
  OR2 C1243 ( .A(n5081), .B(n3916), .Z(n3917) );
  OR2 C1244 ( .A(U162_Z_1), .B(n3917), .Z(n3918) );
  OR2 C1245 ( .A(U162_Z_0), .B(n3918), .Z(n3919) );
  OR2 C1252 ( .A(n4974), .B(n4949), .Z(n3921) );
  OR2 C1253 ( .A(U162_Z_5), .B(n3921), .Z(n3922) );
  OR2 C1254 ( .A(n5020), .B(n3922), .Z(n3923) );
  OR2 C1255 ( .A(n5058), .B(n3923), .Z(n3924) );
  OR2 C1256 ( .A(n5081), .B(n3924), .Z(n3925) );
  OR2 C1257 ( .A(U162_Z_1), .B(n3925), .Z(n3926) );
  OR2 C1258 ( .A(U162_Z_0), .B(n3926), .Z(n3927) );
  OR2 C1267 ( .A(n4974), .B(n4949), .Z(n3929) );
  OR2 C1268 ( .A(n4997), .B(n3929), .Z(n3930) );
  OR2 C1269 ( .A(n5020), .B(n3930), .Z(n3931) );
  OR2 C1270 ( .A(U162_Z_3), .B(n3931), .Z(n3932) );
  OR2 C1271 ( .A(n5081), .B(n3932), .Z(n3933) );
  OR2 C1272 ( .A(n5092), .B(n3933), .Z(n3934) );
  OR2 C1273 ( .A(n5093), .B(n3934), .Z(n3935) );
  OR2 C1277 ( .A(U162_Z_6), .B(U162_Z_7), .Z(n3937) );
  OR2 C1278 ( .A(U162_Z_5), .B(n3937), .Z(n3938) );
  OR2 C1279 ( .A(U162_Z_4), .B(n3938), .Z(n3939) );
  OR2 C1280 ( .A(U162_Z_3), .B(n3939), .Z(n3940) );
  OR2 C1281 ( .A(n5081), .B(n3940), .Z(n3941) );
  OR2 C1282 ( .A(n5092), .B(n3941), .Z(n3942) );
  OR2 C1283 ( .A(U162_Z_0), .B(n3942), .Z(n3943) );
  OR2 C1292 ( .A(n4974), .B(n4949), .Z(n3945) );
  OR2 C1293 ( .A(n4997), .B(n3945), .Z(n3946) );
  OR2 C1294 ( .A(n5020), .B(n3946), .Z(n3947) );
  OR2 C1295 ( .A(n5058), .B(n3947), .Z(n3948) );
  OR2 C1296 ( .A(n5081), .B(n3948), .Z(n3949) );
  OR2 C1297 ( .A(n5092), .B(n3949), .Z(n3950) );
  OR2 C1298 ( .A(U162_Z_0), .B(n3950), .Z(n3951) );
  OR2 C1303 ( .A(U162_Z_14), .B(U162_Z_15), .Z(n3953) );
  OR2 C1304 ( .A(U162_Z_13), .B(n3953), .Z(n3954) );
  OR2 C1305 ( .A(U162_Z_12), .B(n3954), .Z(n3955) );
  OR2 C1306 ( .A(U162_Z_11), .B(n3955), .Z(n3956) );
  OR2 C1307 ( .A(n5091), .B(n3956), .Z(n3957) );
  OR2 C1308 ( .A(n4934), .B(n3957), .Z(n3958) );
  OR2 C1309 ( .A(n4941), .B(n3958), .Z(n3959) );
  OR2 C1316 ( .A(n5087), .B(U162_Z_15), .Z(n3961) );
  OR2 C1317 ( .A(n5088), .B(n3961), .Z(n3962) );
  OR2 C1318 ( .A(n5089), .B(n3962), .Z(n3963) );
  OR2 C1319 ( .A(n5090), .B(n3963), .Z(n3964) );
  OR2 C1320 ( .A(n5091), .B(n3964), .Z(n3965) );
  OR2 C1321 ( .A(U162_Z_9), .B(n3965), .Z(n3966) );
  OR2 C1322 ( .A(U162_Z_8), .B(n3966), .Z(n3967) );
  OR2 C1327 ( .A(U162_Z_14), .B(U162_Z_15), .Z(n3969) );
  OR2 C1328 ( .A(U162_Z_13), .B(n3969), .Z(n3970) );
  OR2 C1329 ( .A(n5089), .B(n3970), .Z(n3971) );
  OR2 C1330 ( .A(n5090), .B(n3971), .Z(n3972) );
  OR2 C1331 ( .A(n5091), .B(n3972), .Z(n3973) );
  OR2 C1332 ( .A(U162_Z_9), .B(n3973), .Z(n3974) );
  OR2 C1333 ( .A(U162_Z_8), .B(n3974), .Z(n3975) );
  OR2 C1340 ( .A(U162_Z_14), .B(n5086), .Z(n3977) );
  OR2 C1341 ( .A(n5088), .B(n3977), .Z(n3978) );
  OR2 C1342 ( .A(n5089), .B(n3978), .Z(n3979) );
  OR2 C1343 ( .A(n5090), .B(n3979), .Z(n3980) );
  OR2 C1344 ( .A(n5091), .B(n3980), .Z(n3981) );
  OR2 C1345 ( .A(U162_Z_9), .B(n3981), .Z(n3982) );
  OR2 C1346 ( .A(U162_Z_8), .B(n3982), .Z(n3983) );
  OR2 C1352 ( .A(U162_Z_14), .B(U162_Z_15), .Z(n3985) );
  OR2 C1353 ( .A(n5088), .B(n3985), .Z(n3986) );
  OR2 C1354 ( .A(n5089), .B(n3986), .Z(n3987) );
  OR2 C1355 ( .A(n5090), .B(n3987), .Z(n3988) );
  OR2 C1356 ( .A(n5091), .B(n3988), .Z(n3989) );
  OR2 C1357 ( .A(U162_Z_9), .B(n3989), .Z(n3990) );
  OR2 C1358 ( .A(U162_Z_8), .B(n3990), .Z(n3991) );
  OR2 C1365 ( .A(n5087), .B(n5086), .Z(n3993) );
  OR2 C1366 ( .A(U162_Z_13), .B(n3993), .Z(n3994) );
  OR2 C1367 ( .A(n5089), .B(n3994), .Z(n3995) );
  OR2 C1368 ( .A(n5090), .B(n3995), .Z(n3996) );
  OR2 C1369 ( .A(n5091), .B(n3996), .Z(n3997) );
  OR2 C1370 ( .A(U162_Z_9), .B(n3997), .Z(n3998) );
  OR2 C1371 ( .A(U162_Z_8), .B(n3998), .Z(n3999) );
  OR2 C1380 ( .A(n5087), .B(n5086), .Z(n4001) );
  OR2 C1381 ( .A(n5088), .B(n4001), .Z(n4002) );
  OR2 C1382 ( .A(n5089), .B(n4002), .Z(n4003) );
  OR2 C1383 ( .A(U162_Z_11), .B(n4003), .Z(n4004) );
  OR2 C1384 ( .A(n5091), .B(n4004), .Z(n4005) );
  OR2 C1385 ( .A(n4934), .B(n4005), .Z(n4006) );
  OR2 C1386 ( .A(n4941), .B(n4006), .Z(n4007) );
  OR2 C1390 ( .A(U162_Z_14), .B(U162_Z_15), .Z(n4009) );
  OR2 C1391 ( .A(U162_Z_13), .B(n4009), .Z(n4010) );
  OR2 C1392 ( .A(U162_Z_12), .B(n4010), .Z(n4011) );
  OR2 C1393 ( .A(U162_Z_11), .B(n4011), .Z(n4012) );
  OR2 C1394 ( .A(n5091), .B(n4012), .Z(n4013) );
  OR2 C1395 ( .A(n4934), .B(n4013), .Z(n4014) );
  OR2 C1396 ( .A(U162_Z_8), .B(n4014), .Z(n4015) );
  OR2 C1405 ( .A(n5087), .B(n5086), .Z(n4017) );
  OR2 C1406 ( .A(n5088), .B(n4017), .Z(n4018) );
  OR2 C1407 ( .A(n5089), .B(n4018), .Z(n4019) );
  OR2 C1408 ( .A(n5090), .B(n4019), .Z(n4020) );
  OR2 C1409 ( .A(n5091), .B(n4020), .Z(n4021) );
  OR2 C1410 ( .A(n4934), .B(n4021), .Z(n4022) );
  OR2 C1411 ( .A(U162_Z_8), .B(n4022), .Z(n4023) );
  OR2 C1416 ( .A(U162_Z_22), .B(U162_Z_23), .Z(n4025) );
  OR2 C1417 ( .A(U162_Z_21), .B(n4025), .Z(n4026) );
  OR2 C1418 ( .A(U162_Z_20), .B(n4026), .Z(n4027) );
  OR2 C1419 ( .A(U162_Z_19), .B(n4027), .Z(n4028) );
  OR2 C1420 ( .A(n5083), .B(n4028), .Z(n4029) );
  OR2 C1421 ( .A(n5084), .B(n4029), .Z(n4030) );
  OR2 C1422 ( .A(n5085), .B(n4030), .Z(n4031) );
  OR2 C1429 ( .A(n5078), .B(U162_Z_23), .Z(n4033) );
  OR2 C1430 ( .A(n5079), .B(n4033), .Z(n4034) );
  OR2 C1431 ( .A(n5080), .B(n4034), .Z(n4035) );
  OR2 C1432 ( .A(n5082), .B(n4035), .Z(n4036) );
  OR2 C1433 ( .A(n5083), .B(n4036), .Z(n4037) );
  OR2 C1434 ( .A(U162_Z_17), .B(n4037), .Z(n4038) );
  OR2 C1435 ( .A(U162_Z_16), .B(n4038), .Z(n4039) );
  OR2 C1440 ( .A(U162_Z_22), .B(U162_Z_23), .Z(n4041) );
  OR2 C1441 ( .A(U162_Z_21), .B(n4041), .Z(n4042) );
  OR2 C1442 ( .A(n5080), .B(n4042), .Z(n4043) );
  OR2 C1443 ( .A(n5082), .B(n4043), .Z(n4044) );
  OR2 C1444 ( .A(n5083), .B(n4044), .Z(n4045) );
  OR2 C1445 ( .A(U162_Z_17), .B(n4045), .Z(n4046) );
  OR2 C1446 ( .A(U162_Z_16), .B(n4046), .Z(n4047) );
  OR2 C1453 ( .A(U162_Z_22), .B(n5070), .Z(n4049) );
  OR2 C1454 ( .A(n5079), .B(n4049), .Z(n4050) );
  OR2 C1455 ( .A(n5080), .B(n4050), .Z(n4051) );
  OR2 C1456 ( .A(n5082), .B(n4051), .Z(n4052) );
  OR2 C1457 ( .A(n5083), .B(n4052), .Z(n4053) );
  OR2 C1458 ( .A(U162_Z_17), .B(n4053), .Z(n4054) );
  OR2 C1459 ( .A(U162_Z_16), .B(n4054), .Z(n4055) );
  OR2 C1465 ( .A(U162_Z_22), .B(U162_Z_23), .Z(n4057) );
  OR2 C1466 ( .A(n5079), .B(n4057), .Z(n4058) );
  OR2 C1467 ( .A(n5080), .B(n4058), .Z(n4059) );
  OR2 C1468 ( .A(n5082), .B(n4059), .Z(n4060) );
  OR2 C1469 ( .A(n5083), .B(n4060), .Z(n4061) );
  OR2 C1470 ( .A(U162_Z_17), .B(n4061), .Z(n4062) );
  OR2 C1471 ( .A(U162_Z_16), .B(n4062), .Z(n4063) );
  OR2 C1478 ( .A(n5078), .B(n5070), .Z(n4065) );
  OR2 C1479 ( .A(U162_Z_21), .B(n4065), .Z(n4066) );
  OR2 C1480 ( .A(n5080), .B(n4066), .Z(n4067) );
  OR2 C1481 ( .A(n5082), .B(n4067), .Z(n4068) );
  OR2 C1482 ( .A(n5083), .B(n4068), .Z(n4069) );
  OR2 C1483 ( .A(U162_Z_17), .B(n4069), .Z(n4070) );
  OR2 C1484 ( .A(U162_Z_16), .B(n4070), .Z(n4071) );
  OR2 C1493 ( .A(n5078), .B(n5070), .Z(n4073) );
  OR2 C1494 ( .A(n5079), .B(n4073), .Z(n4074) );
  OR2 C1495 ( .A(n5080), .B(n4074), .Z(n4075) );
  OR2 C1496 ( .A(U162_Z_19), .B(n4075), .Z(n4076) );
  OR2 C1497 ( .A(n5083), .B(n4076), .Z(n4077) );
  OR2 C1498 ( .A(n5084), .B(n4077), .Z(n4078) );
  OR2 C1499 ( .A(n5085), .B(n4078), .Z(n4079) );
  OR2 C1503 ( .A(U162_Z_22), .B(U162_Z_23), .Z(n4081) );
  OR2 C1504 ( .A(U162_Z_21), .B(n4081), .Z(n4082) );
  OR2 C1505 ( .A(U162_Z_20), .B(n4082), .Z(n4083) );
  OR2 C1506 ( .A(U162_Z_19), .B(n4083), .Z(n4084) );
  OR2 C1507 ( .A(n5083), .B(n4084), .Z(n4085) );
  OR2 C1508 ( .A(n5084), .B(n4085), .Z(n4086) );
  OR2 C1509 ( .A(U162_Z_16), .B(n4086), .Z(n4087) );
  OR2 C1518 ( .A(n5078), .B(n5070), .Z(n4089) );
  OR2 C1519 ( .A(n5079), .B(n4089), .Z(n4090) );
  OR2 C1520 ( .A(n5080), .B(n4090), .Z(n4091) );
  OR2 C1521 ( .A(n5082), .B(n4091), .Z(n4092) );
  OR2 C1522 ( .A(n5083), .B(n4092), .Z(n4093) );
  OR2 C1523 ( .A(n5084), .B(n4093), .Z(n4094) );
  OR2 C1524 ( .A(U162_Z_16), .B(n4094), .Z(n4095) );
  OR2 C1529 ( .A(U162_Z_30), .B(U162_Z_31), .Z(n4097) );
  OR2 C1530 ( .A(U162_Z_29), .B(n4097), .Z(n4098) );
  OR2 C1531 ( .A(U162_Z_28), .B(n4098), .Z(n4099) );
  OR2 C1532 ( .A(U162_Z_27), .B(n4099), .Z(n4100) );
  OR2 C1533 ( .A(n5062), .B(n4100), .Z(n4101) );
  OR2 C1534 ( .A(n5063), .B(n4101), .Z(n4102) );
  OR2 C1535 ( .A(n5064), .B(n4102), .Z(n4103) );
  OR2 C1542 ( .A(n5057), .B(U162_Z_31), .Z(n4105) );
  OR2 C1543 ( .A(n5059), .B(n4105), .Z(n4106) );
  OR2 C1544 ( .A(n5060), .B(n4106), .Z(n4107) );
  OR2 C1545 ( .A(n5061), .B(n4107), .Z(n4108) );
  OR2 C1546 ( .A(n5062), .B(n4108), .Z(n4109) );
  OR2 C1547 ( .A(U162_Z_25), .B(n4109), .Z(n4110) );
  OR2 C1548 ( .A(U162_Z_24), .B(n4110), .Z(n4111) );
  OR2 C1553 ( .A(U162_Z_30), .B(U162_Z_31), .Z(n4113) );
  OR2 C1554 ( .A(U162_Z_29), .B(n4113), .Z(n4114) );
  OR2 C1555 ( .A(n5060), .B(n4114), .Z(n4115) );
  OR2 C1556 ( .A(n5061), .B(n4115), .Z(n4116) );
  OR2 C1557 ( .A(n5062), .B(n4116), .Z(n4117) );
  OR2 C1558 ( .A(U162_Z_25), .B(n4117), .Z(n4118) );
  OR2 C1559 ( .A(U162_Z_24), .B(n4118), .Z(n4119) );
  OR2 C1566 ( .A(U162_Z_30), .B(n5049), .Z(n4121) );
  OR2 C1567 ( .A(n5059), .B(n4121), .Z(n4122) );
  OR2 C1568 ( .A(n5060), .B(n4122), .Z(n4123) );
  OR2 C1569 ( .A(n5061), .B(n4123), .Z(n4124) );
  OR2 C1570 ( .A(n5062), .B(n4124), .Z(n4125) );
  OR2 C1571 ( .A(U162_Z_25), .B(n4125), .Z(n4126) );
  OR2 C1572 ( .A(U162_Z_24), .B(n4126), .Z(n4127) );
  OR2 C1578 ( .A(U162_Z_30), .B(U162_Z_31), .Z(n4129) );
  OR2 C1579 ( .A(n5059), .B(n4129), .Z(n4130) );
  OR2 C1580 ( .A(n5060), .B(n4130), .Z(n4131) );
  OR2 C1581 ( .A(n5061), .B(n4131), .Z(n4132) );
  OR2 C1582 ( .A(n5062), .B(n4132), .Z(n4133) );
  OR2 C1583 ( .A(U162_Z_25), .B(n4133), .Z(n4134) );
  OR2 C1584 ( .A(U162_Z_24), .B(n4134), .Z(n4135) );
  OR2 C1591 ( .A(n5057), .B(n5049), .Z(n4137) );
  OR2 C1592 ( .A(U162_Z_29), .B(n4137), .Z(n4138) );
  OR2 C1593 ( .A(n5060), .B(n4138), .Z(n4139) );
  OR2 C1594 ( .A(n5061), .B(n4139), .Z(n4140) );
  OR2 C1595 ( .A(n5062), .B(n4140), .Z(n4141) );
  OR2 C1596 ( .A(U162_Z_25), .B(n4141), .Z(n4142) );
  OR2 C1597 ( .A(U162_Z_24), .B(n4142), .Z(n4143) );
  OR2 C1606 ( .A(n5057), .B(n5049), .Z(n4145) );
  OR2 C1607 ( .A(n5059), .B(n4145), .Z(n4146) );
  OR2 C1608 ( .A(n5060), .B(n4146), .Z(n4147) );
  OR2 C1609 ( .A(U162_Z_27), .B(n4147), .Z(n4148) );
  OR2 C1610 ( .A(n5062), .B(n4148), .Z(n4149) );
  OR2 C1611 ( .A(n5063), .B(n4149), .Z(n4150) );
  OR2 C1612 ( .A(n5064), .B(n4150), .Z(n4151) );
  OR2 C1616 ( .A(U162_Z_30), .B(U162_Z_31), .Z(n4153) );
  OR2 C1617 ( .A(U162_Z_29), .B(n4153), .Z(n4154) );
  OR2 C1618 ( .A(U162_Z_28), .B(n4154), .Z(n4155) );
  OR2 C1619 ( .A(U162_Z_27), .B(n4155), .Z(n4156) );
  OR2 C1620 ( .A(n5062), .B(n4156), .Z(n4157) );
  OR2 C1621 ( .A(n5063), .B(n4157), .Z(n4158) );
  OR2 C1622 ( .A(U162_Z_24), .B(n4158), .Z(n4159) );
  OR2 C1631 ( .A(n5057), .B(n5049), .Z(n4161) );
  OR2 C1632 ( .A(n5059), .B(n4161), .Z(n4162) );
  OR2 C1633 ( .A(n5060), .B(n4162), .Z(n4163) );
  OR2 C1634 ( .A(n5061), .B(n4163), .Z(n4164) );
  OR2 C1635 ( .A(n5062), .B(n4164), .Z(n4165) );
  OR2 C1636 ( .A(n5063), .B(n4165), .Z(n4166) );
  OR2 C1637 ( .A(U162_Z_24), .B(n4166), .Z(n4167) );
  OR2 C1649 ( .A(n5457), .B(U157_CONTROL2), .Z(n4170) );
  OR2 C1687 ( .A(n5458), .B(n5457), .Z(n4172) );
  OR2 C1767 ( .A(n3267), .B(n3268), .Z(n4173) );
  IV I_196 ( .A(reset_to_pma_tx), .Z(n3179) );
  AN2 C1828 ( .A(U161_Z_0), .B(n4948), .Z(n3197) );
  AN2 C1829 ( .A(U161_Z_1), .B(n4940), .Z(n3198) );
  AN2 C1830 ( .A(U161_Z_2), .B(n5069), .Z(n3199) );
  AN2 C1831 ( .A(U161_Z_3), .B(n5048), .Z(n3200) );
  AN2 C1832 ( .A(U161_Z_4), .B(n5027), .Z(n3201) );
  AN2 C1833 ( .A(U161_Z_5), .B(n5004), .Z(n3202) );
  AN2 C1834 ( .A(U161_Z_6), .B(n4983), .Z(n3203) );
  AN2 C1835 ( .A(U161_Z_7), .B(n4962), .Z(n3204) );
  AN2 C1836 ( .A(n5102), .B(n4175), .Z(n3205) );
  OR2 C1837 ( .A(n4946), .B(n4957), .Z(n4175) );
  AN2 C1838 ( .A(n5095), .B(n4176), .Z(n3206) );
  OR2 C1839 ( .A(n5025), .B(n5036), .Z(n4176) );
  AN2 C1840 ( .A(n5097), .B(n4947), .Z(n3207) );
  AN2 C1841 ( .A(n5096), .B(n5026), .Z(n3208) );
  AN2 C1842 ( .A(U161_Z_0), .B(n4942), .Z(n3209) );
  AN2 C1843 ( .A(U161_Z_1), .B(n4924), .Z(n3210) );
  AN2 C1844 ( .A(U161_Z_2), .B(n5065), .Z(n3211) );
  AN2 C1845 ( .A(U161_Z_3), .B(n5044), .Z(n3212) );
  AN2 C1846 ( .A(U161_Z_4), .B(n5021), .Z(n3213) );
  AN2 C1847 ( .A(U161_Z_5), .B(n5000), .Z(n3214) );
  AN2 C1848 ( .A(U161_Z_6), .B(n4979), .Z(n3215) );
  AN2 C1849 ( .A(U161_Z_7), .B(n4958), .Z(n3216) );
  AN2 C1850 ( .A(U161_Z_0), .B(n4956), .Z(n3224) );
  AN2 C1851 ( .A(U161_Z_1), .B(n4933), .Z(n3223) );
  AN2 C1852 ( .A(U161_Z_2), .B(n5077), .Z(n3222) );
  AN2 C1853 ( .A(U161_Z_3), .B(n5056), .Z(n3221) );
  AN2 C1854 ( .A(U161_Z_4), .B(n5035), .Z(n3220) );
  AN2 C1855 ( .A(U161_Z_5), .B(n5012), .Z(n3219) );
  AN2 C1856 ( .A(U161_Z_6), .B(n4991), .Z(n3218) );
  AN2 C1857 ( .A(U161_Z_7), .B(n4970), .Z(n3217) );
  AN2 C1858 ( .A(U161_Z_0), .B(n4183), .Z(n3225) );
  OR2 C1859 ( .A(n4182), .B(n4950), .Z(n4183) );
  OR2 C1860 ( .A(n4181), .B(n4943), .Z(n4182) );
  OR2 C1861 ( .A(n4180), .B(n4944), .Z(n4181) );
  OR2 C1862 ( .A(n4179), .B(n4951), .Z(n4180) );
  OR2 C1863 ( .A(n4178), .B(n4945), .Z(n4179) );
  OR2 C1864 ( .A(n4177), .B(n4952), .Z(n4178) );
  OR2 C1865 ( .A(n4954), .B(n4953), .Z(n4177) );
  AN2 C1866 ( .A(U161_Z_1), .B(n4190), .Z(n3226) );
  OR2 C1867 ( .A(n4189), .B(n4925), .Z(n4190) );
  OR2 C1868 ( .A(n4188), .B(n4926), .Z(n4189) );
  OR2 C1869 ( .A(n4187), .B(n4935), .Z(n4188) );
  OR2 C1870 ( .A(n4186), .B(n4936), .Z(n4187) );
  OR2 C1871 ( .A(n4185), .B(n4937), .Z(n4186) );
  OR2 C1872 ( .A(n4184), .B(n4938), .Z(n4185) );
  OR2 C1873 ( .A(n4927), .B(n4939), .Z(n4184) );
  AN2 C1874 ( .A(U161_Z_2), .B(n4197), .Z(n3227) );
  OR2 C1875 ( .A(n4196), .B(n5071), .Z(n4197) );
  OR2 C1876 ( .A(n4195), .B(n5066), .Z(n4196) );
  OR2 C1877 ( .A(n4194), .B(n5067), .Z(n4195) );
  OR2 C1878 ( .A(n4193), .B(n5072), .Z(n4194) );
  OR2 C1879 ( .A(n4192), .B(n5068), .Z(n4193) );
  OR2 C1880 ( .A(n4191), .B(n5073), .Z(n4192) );
  OR2 C1881 ( .A(n5075), .B(n5074), .Z(n4191) );
  AN2 C1882 ( .A(U161_Z_3), .B(n4204), .Z(n3228) );
  OR2 C1883 ( .A(n4203), .B(n5050), .Z(n4204) );
  OR2 C1884 ( .A(n4202), .B(n5045), .Z(n4203) );
  OR2 C1885 ( .A(n4201), .B(n5046), .Z(n4202) );
  OR2 C1886 ( .A(n4200), .B(n5051), .Z(n4201) );
  OR2 C1887 ( .A(n4199), .B(n5047), .Z(n4200) );
  OR2 C1888 ( .A(n4198), .B(n5052), .Z(n4199) );
  OR2 C1889 ( .A(n5054), .B(n5053), .Z(n4198) );
  AN2 C1890 ( .A(U161_Z_4), .B(n4211), .Z(n3229) );
  OR2 C1891 ( .A(n4210), .B(n5029), .Z(n4211) );
  OR2 C1892 ( .A(n4209), .B(n5022), .Z(n4210) );
  OR2 C1893 ( .A(n4208), .B(n5023), .Z(n4209) );
  OR2 C1894 ( .A(n4207), .B(n5030), .Z(n4208) );
  OR2 C1895 ( .A(n4206), .B(n5024), .Z(n4207) );
  OR2 C1896 ( .A(n4205), .B(n5031), .Z(n4206) );
  OR2 C1897 ( .A(n5033), .B(n5032), .Z(n4205) );
  AN2 C1898 ( .A(U161_Z_5), .B(n4218), .Z(n3230) );
  OR2 C1899 ( .A(n4217), .B(n5006), .Z(n4218) );
  OR2 C1900 ( .A(n4216), .B(n5001), .Z(n4217) );
  OR2 C1901 ( .A(n4215), .B(n5002), .Z(n4216) );
  OR2 C1902 ( .A(n4214), .B(n5007), .Z(n4215) );
  OR2 C1903 ( .A(n4213), .B(n5003), .Z(n4214) );
  OR2 C1904 ( .A(n4212), .B(n5008), .Z(n4213) );
  OR2 C1905 ( .A(n5010), .B(n5009), .Z(n4212) );
  AN2 C1906 ( .A(U161_Z_6), .B(n4225), .Z(n3231) );
  OR2 C1907 ( .A(n4224), .B(n4985), .Z(n4225) );
  OR2 C1908 ( .A(n4223), .B(n4980), .Z(n4224) );
  OR2 C1909 ( .A(n4222), .B(n4981), .Z(n4223) );
  OR2 C1910 ( .A(n4221), .B(n4986), .Z(n4222) );
  OR2 C1911 ( .A(n4220), .B(n4982), .Z(n4221) );
  OR2 C1912 ( .A(n4219), .B(n4987), .Z(n4220) );
  OR2 C1913 ( .A(n4989), .B(n4988), .Z(n4219) );
  AN2 C1914 ( .A(U161_Z_7), .B(n4232), .Z(n3232) );
  OR2 C1915 ( .A(n4231), .B(n4964), .Z(n4232) );
  OR2 C1916 ( .A(n4230), .B(n4959), .Z(n4231) );
  OR2 C1917 ( .A(n4229), .B(n4960), .Z(n4230) );
  OR2 C1918 ( .A(n4228), .B(n4965), .Z(n4229) );
  OR2 C1919 ( .A(n4227), .B(n4961), .Z(n4228) );
  OR2 C1920 ( .A(n4226), .B(n4966), .Z(n4227) );
  OR2 C1921 ( .A(n4968), .B(n4967), .Z(n4226) );
  OR2 C1922 ( .A(n3225), .B(n3209), .Z(n3233) );
  OR2 C1923 ( .A(n3226), .B(n3210), .Z(n3234) );
  OR2 C1924 ( .A(n3227), .B(n3211), .Z(n3235) );
  OR2 C1925 ( .A(n3228), .B(n3212), .Z(n3236) );
  OR2 C1926 ( .A(n3229), .B(n3213), .Z(n3237) );
  OR2 C1927 ( .A(n3230), .B(n3214), .Z(n3238) );
  OR2 C1928 ( .A(n3231), .B(n3215), .Z(n3239) );
  OR2 C1929 ( .A(n3232), .B(n3216), .Z(n3240) );
  AN2 C1930 ( .A(n5105), .B(n5104), .Z(n3241) );
  AN2 C1931 ( .A(n3241), .B(n5103), .Z(n3242) );
  AN2 C1932 ( .A(n3242), .B(n3200), .Z(n3243) );
  AN2 C1933 ( .A(n3242), .B(n5101), .Z(n3244) );
  AN2 C1934 ( .A(n3244), .B(n5100), .Z(n3245) );
  AN2 C1935 ( .A(n3245), .B(n5099), .Z(n3246) );
  AN2 C1936 ( .A(n3246), .B(n5098), .Z(n3247) );
  AN2 C1937 ( .A(n3476), .B(n5453), .Z(n3248) );
  OR2 C1939 ( .A(n4252), .B(n4253), .Z(n3249) );
  OR2 C1940 ( .A(n4247), .B(n4251), .Z(n4252) );
  OR2 C1941 ( .A(n4242), .B(n4246), .Z(n4247) );
  AN2 C1942 ( .A(n4239), .B(n4241), .Z(n4242) );
  AN2 C1943 ( .A(n4238), .B(n3232), .Z(n4239) );
  AN2 C1944 ( .A(n4237), .B(n3231), .Z(n4238) );
  AN2 C1945 ( .A(n4236), .B(n3230), .Z(n4237) );
  AN2 C1946 ( .A(n4235), .B(n3229), .Z(n4236) );
  AN2 C1947 ( .A(n4234), .B(n3228), .Z(n4235) );
  AN2 C1948 ( .A(n4233), .B(n3227), .Z(n4234) );
  AN2 C1949 ( .A(n3225), .B(n3226), .Z(n4233) );
  OR2 C1950 ( .A(n4240), .B(n4928), .Z(n4241) );
  OR2 C1951 ( .A(n4932), .B(n4931), .Z(n4240) );
  AN2 C1952 ( .A(n4245), .B(n3240), .Z(n4246) );
  AN2 C1953 ( .A(n4244), .B(n3239), .Z(n4245) );
  AN2 C1954 ( .A(n4243), .B(n3238), .Z(n4244) );
  AN2 C1955 ( .A(n3205), .B(n3237), .Z(n4243) );
  AN2 C1956 ( .A(n4250), .B(n3236), .Z(n4251) );
  AN2 C1957 ( .A(n4249), .B(n3235), .Z(n4250) );
  AN2 C1958 ( .A(n4248), .B(n3234), .Z(n4249) );
  AN2 C1959 ( .A(n3206), .B(n3233), .Z(n4248) );
  AN2 C1960 ( .A(n3205), .B(n3206), .Z(n4253) );
  AN2 C1961 ( .A(n4259), .B(n3217), .Z(n3250) );
  AN2 C1962 ( .A(n4258), .B(n3218), .Z(n4259) );
  AN2 C1963 ( .A(n4257), .B(n3219), .Z(n4258) );
  AN2 C1964 ( .A(n4256), .B(n3220), .Z(n4257) );
  AN2 C1965 ( .A(n4255), .B(n3221), .Z(n4256) );
  AN2 C1966 ( .A(n4254), .B(n3222), .Z(n4255) );
  AN2 C1967 ( .A(n3224), .B(n3223), .Z(n4254) );
  OR2 C1968 ( .A(n3207), .B(n4264), .Z(n3251) );
  AN2 C1969 ( .A(n3208), .B(n4263), .Z(n4264) );
  OR2 C1970 ( .A(n3205), .B(n4262), .Z(n4263) );
  AN2 C1971 ( .A(n4261), .B(n3236), .Z(n4262) );
  AN2 C1972 ( .A(n4260), .B(n3235), .Z(n4261) );
  AN2 C1973 ( .A(n3233), .B(n3234), .Z(n4260) );
  OR2 C1974 ( .A(n4311), .B(n4312), .Z(n3252) );
  OR2 C1975 ( .A(n4308), .B(n4310), .Z(n4311) );
  OR2 C1976 ( .A(n4304), .B(n4307), .Z(n4308) );
  OR2 C1977 ( .A(n4299), .B(n4303), .Z(n4304) );
  OR2 C1978 ( .A(n4293), .B(n4298), .Z(n4299) );
  OR2 C1979 ( .A(n4286), .B(n4292), .Z(n4293) );
  OR2 C1980 ( .A(n4279), .B(n4285), .Z(n4286) );
  OR2 C1981 ( .A(n4271), .B(n4278), .Z(n4279) );
  AN2 C1982 ( .A(n4270), .B(n3240), .Z(n4271) );
  AN2 C1983 ( .A(n4269), .B(n3239), .Z(n4270) );
  AN2 C1984 ( .A(n4268), .B(n3238), .Z(n4269) );
  AN2 C1985 ( .A(n4267), .B(n3237), .Z(n4268) );
  AN2 C1986 ( .A(n4266), .B(n3236), .Z(n4267) );
  AN2 C1987 ( .A(n4265), .B(n3235), .Z(n4266) );
  AN2 C1988 ( .A(n3197), .B(n3234), .Z(n4265) );
  AN2 C1989 ( .A(n4277), .B(n3240), .Z(n4278) );
  AN2 C1990 ( .A(n4276), .B(n3239), .Z(n4277) );
  AN2 C1991 ( .A(n4275), .B(n3238), .Z(n4276) );
  AN2 C1992 ( .A(n4274), .B(n3237), .Z(n4275) );
  AN2 C1993 ( .A(n4273), .B(n3236), .Z(n4274) );
  AN2 C1994 ( .A(n4272), .B(n3235), .Z(n4273) );
  AN2 C1995 ( .A(n5105), .B(n3198), .Z(n4272) );
  AN2 C1996 ( .A(n4284), .B(n3240), .Z(n4285) );
  AN2 C1997 ( .A(n4283), .B(n3239), .Z(n4284) );
  AN2 C1998 ( .A(n4282), .B(n3238), .Z(n4283) );
  AN2 C1999 ( .A(n4281), .B(n3237), .Z(n4282) );
  AN2 C2000 ( .A(n4280), .B(n3236), .Z(n4281) );
  AN2 C2001 ( .A(n3241), .B(n3199), .Z(n4280) );
  AN2 C2002 ( .A(n4290), .B(n4291), .Z(n4292) );
  AN2 C2003 ( .A(n4289), .B(n3240), .Z(n4290) );
  AN2 C2004 ( .A(n4288), .B(n3239), .Z(n4289) );
  AN2 C2005 ( .A(n4287), .B(n3238), .Z(n4288) );
  AN2 C2006 ( .A(n3243), .B(n3237), .Z(n4287) );
  IV I_205 ( .A(ALTERNATE_ENCODE), .Z(n4291) );
  AN2 C2008 ( .A(n4297), .B(ALTERNATE_ENCODE), .Z(n4298) );
  AN2 C2009 ( .A(n4296), .B(n5094), .Z(n4297) );
  AN2 C2010 ( .A(n4295), .B(n5098), .Z(n4296) );
  AN2 C2011 ( .A(n4294), .B(n5099), .Z(n4295) );
  AN2 C2012 ( .A(n3243), .B(n3206), .Z(n4294) );
  AN2 C2013 ( .A(n4302), .B(n3240), .Z(n4303) );
  AN2 C2014 ( .A(n4301), .B(n3239), .Z(n4302) );
  AN2 C2015 ( .A(n4300), .B(n3238), .Z(n4301) );
  AN2 C2016 ( .A(n3244), .B(n3201), .Z(n4300) );
  AN2 C2017 ( .A(n4306), .B(n3240), .Z(n4307) );
  AN2 C2018 ( .A(n4305), .B(n3239), .Z(n4306) );
  AN2 C2019 ( .A(n3245), .B(n3202), .Z(n4305) );
  AN2 C2020 ( .A(n4309), .B(n3240), .Z(n4310) );
  AN2 C2021 ( .A(n3246), .B(n3203), .Z(n4309) );
  AN2 C2022 ( .A(n3247), .B(n3204), .Z(n4312) );
  AN2 C2023 ( .A(n3247), .B(n5094), .Z(n3253) );
  AN2 C218 ( .A(n4396), .B(n4395), .Z(n4366) );
  AN2 C217 ( .A(n4366), .B(n4394), .Z(n4365) );
  AN2 C216 ( .A(n4365), .B(n4393), .Z(n4364) );
  AN2 C215 ( .A(n4364), .B(n4392), .Z(n4363) );
  AN2 C214 ( .A(n4363), .B(n4391), .Z(n4362) );
  AN2 C213 ( .A(n4362), .B(n4390), .Z(n4361) );
  AN2 C212 ( .A(n4361), .B(n4389), .Z(n4360) );
  AN2 C211 ( .A(n4360), .B(n4388), .Z(n4359) );
  AN2 C210 ( .A(n4359), .B(n4387), .Z(n4358) );
  AN2 C209 ( .A(n4358), .B(n4379), .Z(n4357) );
  AN2 C208 ( .A(n4357), .B(n5275), .Z(n4356) );
  AN2 C207 ( .A(n4356), .B(tx_fifo_pop_pre), .Z(assertion_shengyushen) );
  OR2 C206 ( .A(loopback_xgmii), .B(n4476), .Z(n4367) );
  OR2 C205 ( .A(n4367), .B(reset_to_xgmii_tx), .Z(n4398) );
  AN2 C204 ( .A(tx_test_pat_en), .B(test_pat_sel), .Z(n4476) );
  AN2 C202 ( .A(tx_test_pat_en), .B(n4393), .Z(n4477) );
  OR2 C199 ( .A(n4480), .B(n5476), .Z(n4479) );
  OR2 C190 ( .A(tx_mode[0]), .B(n5477), .Z(n4369) );
  OR2 C187 ( .A(U155_Z_0), .B(n4373), .Z(n4372) );
  OR2 C186 ( .A(U154_Z_0), .B(n4374), .Z(n4373) );
  OR2 C185 ( .A(U154_Z_1), .B(n4375), .Z(n4374) );
  OR2 C184 ( .A(U154_Z_2), .B(n4376), .Z(n4375) );
  OR2 C183 ( .A(U155_Z_1), .B(n4377), .Z(n4376) );
  OR2 C182 ( .A(U154_Z_3), .B(n4378), .Z(n4377) );
  OR2 C181 ( .A(U154_Z_4), .B(U154_Z_5), .Z(n4378) );
  IV I_10 ( .A(n4380), .Z(n4379) );
  OR2 C179 ( .A(txc_xfi[0]), .B(n4381), .Z(n4380) );
  OR2 C178 ( .A(txc_xfi[1]), .B(n4382), .Z(n4381) );
  OR2 C177 ( .A(txc_xfi[2]), .B(n4383), .Z(n4382) );
  OR2 C176 ( .A(txc_xfi[3]), .B(n4384), .Z(n4383) );
  OR2 C175 ( .A(txc_xfi[4]), .B(n4385), .Z(n4384) );
  OR2 C174 ( .A(txc_xfi[5]), .B(n4386), .Z(n4385) );
  OR2 C173 ( .A(txc_xfi[6]), .B(txc_xfi[7]), .Z(n4386) );
  IV I_9 ( .A(ALTERNATE_ENCODE), .Z(n4387) );
  IV I_8 ( .A(scr_bypass_enable), .Z(n4388) );
  IV I_7 ( .A(data_pat_sel), .Z(n4389) );
  IV I_6 ( .A(tx_prbs_pat_en), .Z(n4390) );
  IV I_5 ( .A(reset_to_pma_tx), .Z(n4391) );
  IV I_4 ( .A(reset_to_xgmii_tx), .Z(n4392) );
  IV I_3 ( .A(test_pat_sel), .Z(n4393) );
  IV I_2 ( .A(loopback_xgmii), .Z(n4394) );
  IV I_1 ( .A(tx_test_pat_en), .Z(n4395) );
  IV I_0 ( .A(enable_alternate_refresh), .Z(n4396) );
  FD1 test_mode_enc_reg ( .D(n4477), .CP(pma_tx_clk), .Q(n4399) );
  FD1 square_wave_reg ( .D(n4398), .CP(pma_tx_clk), .Q(n4397) );
  FD1 cntl_xfi_reg_0_ ( .D(U161_Z_0), .CP(pma_tx_clk), .Q(U161_DATA3_0) );
  FD1 cntl_xfi_reg_1_ ( .D(U161_Z_1), .CP(pma_tx_clk), .Q(U161_DATA3_1) );
  FD1 cntl_xfi_reg_2_ ( .D(U161_Z_2), .CP(pma_tx_clk), .Q(U161_DATA3_2) );
  FD1 cntl_xfi_reg_3_ ( .D(U161_Z_3), .CP(pma_tx_clk), .Q(U161_DATA3_3) );
  FD1 cntl_xfi_reg_4_ ( .D(U161_Z_4), .CP(pma_tx_clk), .Q(U161_DATA3_4) );
  FD1 cntl_xfi_reg_5_ ( .D(U161_Z_5), .CP(pma_tx_clk), .Q(U161_DATA3_5) );
  FD1 cntl_xfi_reg_6_ ( .D(U161_Z_6), .CP(pma_tx_clk), .Q(U161_DATA3_6) );
  FD1 cntl_xfi_reg_7_ ( .D(U161_Z_7), .CP(pma_tx_clk), .Q(U161_DATA3_7) );
  FD1 data_xfi_reg_0_ ( .D(U162_Z_0), .CP(pma_tx_clk), .Q(U162_DATA3_0) );
  FD1 data_xfi_reg_1_ ( .D(U162_Z_1), .CP(pma_tx_clk), .Q(U162_DATA3_1) );
  FD1 data_xfi_reg_2_ ( .D(U162_Z_2), .CP(pma_tx_clk), .Q(U162_DATA3_2) );
  FD1 data_xfi_reg_3_ ( .D(U162_Z_3), .CP(pma_tx_clk), .Q(U162_DATA3_3) );
  FD1 data_xfi_reg_4_ ( .D(U162_Z_4), .CP(pma_tx_clk), .Q(U162_DATA3_4) );
  FD1 data_xfi_reg_5_ ( .D(U162_Z_5), .CP(pma_tx_clk), .Q(U162_DATA3_5) );
  FD1 data_xfi_reg_6_ ( .D(U162_Z_6), .CP(pma_tx_clk), .Q(U162_DATA3_6) );
  FD1 data_xfi_reg_7_ ( .D(U162_Z_7), .CP(pma_tx_clk), .Q(U162_DATA3_7) );
  FD1 data_xfi_reg_8_ ( .D(U162_Z_8), .CP(pma_tx_clk), .Q(U162_DATA3_8) );
  FD1 data_xfi_reg_9_ ( .D(U162_Z_9), .CP(pma_tx_clk), .Q(U162_DATA3_9) );
  FD1 data_xfi_reg_10_ ( .D(U162_Z_10), .CP(pma_tx_clk), .Q(U162_DATA3_10) );
  FD1 data_xfi_reg_11_ ( .D(U162_Z_11), .CP(pma_tx_clk), .Q(U162_DATA3_11) );
  FD1 data_xfi_reg_12_ ( .D(U162_Z_12), .CP(pma_tx_clk), .Q(U162_DATA3_12) );
  FD1 data_xfi_reg_13_ ( .D(U162_Z_13), .CP(pma_tx_clk), .Q(U162_DATA3_13) );
  FD1 data_xfi_reg_14_ ( .D(U162_Z_14), .CP(pma_tx_clk), .Q(U162_DATA3_14) );
  FD1 data_xfi_reg_15_ ( .D(U162_Z_15), .CP(pma_tx_clk), .Q(U162_DATA3_15) );
  FD1 data_xfi_reg_16_ ( .D(U162_Z_16), .CP(pma_tx_clk), .Q(U162_DATA3_16) );
  FD1 data_xfi_reg_17_ ( .D(U162_Z_17), .CP(pma_tx_clk), .Q(U162_DATA3_17) );
  FD1 data_xfi_reg_18_ ( .D(U162_Z_18), .CP(pma_tx_clk), .Q(U162_DATA3_18) );
  FD1 data_xfi_reg_19_ ( .D(U162_Z_19), .CP(pma_tx_clk), .Q(U162_DATA3_19) );
  FD1 data_xfi_reg_20_ ( .D(U162_Z_20), .CP(pma_tx_clk), .Q(U162_DATA3_20) );
  FD1 data_xfi_reg_21_ ( .D(U162_Z_21), .CP(pma_tx_clk), .Q(U162_DATA3_21) );
  FD1 data_xfi_reg_22_ ( .D(U162_Z_22), .CP(pma_tx_clk), .Q(U162_DATA3_22) );
  FD1 data_xfi_reg_23_ ( .D(U162_Z_23), .CP(pma_tx_clk), .Q(U162_DATA3_23) );
  FD1 data_xfi_reg_24_ ( .D(U162_Z_24), .CP(pma_tx_clk), .Q(U162_DATA3_24) );
  FD1 data_xfi_reg_25_ ( .D(U162_Z_25), .CP(pma_tx_clk), .Q(U162_DATA3_25) );
  FD1 data_xfi_reg_26_ ( .D(U162_Z_26), .CP(pma_tx_clk), .Q(U162_DATA3_26) );
  FD1 data_xfi_reg_27_ ( .D(U162_Z_27), .CP(pma_tx_clk), .Q(U162_DATA3_27) );
  FD1 data_xfi_reg_28_ ( .D(U162_Z_28), .CP(pma_tx_clk), .Q(U162_DATA3_28) );
  FD1 data_xfi_reg_29_ ( .D(U162_Z_29), .CP(pma_tx_clk), .Q(U162_DATA3_29) );
  FD1 data_xfi_reg_30_ ( .D(U162_Z_30), .CP(pma_tx_clk), .Q(U162_DATA3_30) );
  FD1 data_xfi_reg_31_ ( .D(U162_Z_31), .CP(pma_tx_clk), .Q(U162_DATA3_31) );
  FD1 data_xfi_reg_32_ ( .D(U162_Z_32), .CP(pma_tx_clk), .Q(U162_DATA3_32) );
  FD1 data_xfi_reg_33_ ( .D(U162_Z_33), .CP(pma_tx_clk), .Q(U162_DATA3_33) );
  FD1 data_xfi_reg_34_ ( .D(U162_Z_34), .CP(pma_tx_clk), .Q(U162_DATA3_34) );
  FD1 data_xfi_reg_35_ ( .D(U162_Z_35), .CP(pma_tx_clk), .Q(U162_DATA3_35) );
  FD1 data_xfi_reg_36_ ( .D(U162_Z_36), .CP(pma_tx_clk), .Q(U162_DATA3_36) );
  FD1 data_xfi_reg_37_ ( .D(U162_Z_37), .CP(pma_tx_clk), .Q(U162_DATA3_37) );
  FD1 data_xfi_reg_38_ ( .D(U162_Z_38), .CP(pma_tx_clk), .Q(U162_DATA3_38) );
  FD1 data_xfi_reg_39_ ( .D(U162_Z_39), .CP(pma_tx_clk), .Q(U162_DATA3_39) );
  FD1 data_xfi_reg_40_ ( .D(U162_Z_40), .CP(pma_tx_clk), .Q(U162_DATA3_40) );
  FD1 data_xfi_reg_41_ ( .D(U162_Z_41), .CP(pma_tx_clk), .Q(U162_DATA3_41) );
  FD1 data_xfi_reg_42_ ( .D(U162_Z_42), .CP(pma_tx_clk), .Q(U162_DATA3_42) );
  FD1 data_xfi_reg_43_ ( .D(U162_Z_43), .CP(pma_tx_clk), .Q(U162_DATA3_43) );
  FD1 data_xfi_reg_44_ ( .D(U162_Z_44), .CP(pma_tx_clk), .Q(U162_DATA3_44) );
  FD1 data_xfi_reg_45_ ( .D(U162_Z_45), .CP(pma_tx_clk), .Q(U162_DATA3_45) );
  FD1 data_xfi_reg_46_ ( .D(U162_Z_46), .CP(pma_tx_clk), .Q(U162_DATA3_46) );
  FD1 data_xfi_reg_47_ ( .D(U162_Z_47), .CP(pma_tx_clk), .Q(U162_DATA3_47) );
  FD1 data_xfi_reg_48_ ( .D(U162_Z_48), .CP(pma_tx_clk), .Q(U162_DATA3_48) );
  FD1 data_xfi_reg_49_ ( .D(U162_Z_49), .CP(pma_tx_clk), .Q(U162_DATA3_49) );
  FD1 data_xfi_reg_50_ ( .D(U162_Z_50), .CP(pma_tx_clk), .Q(U162_DATA3_50) );
  FD1 data_xfi_reg_51_ ( .D(U162_Z_51), .CP(pma_tx_clk), .Q(U162_DATA3_51) );
  FD1 data_xfi_reg_52_ ( .D(U162_Z_52), .CP(pma_tx_clk), .Q(U162_DATA3_52) );
  FD1 data_xfi_reg_53_ ( .D(U162_Z_53), .CP(pma_tx_clk), .Q(U162_DATA3_53) );
  FD1 data_xfi_reg_54_ ( .D(U162_Z_54), .CP(pma_tx_clk), .Q(U162_DATA3_54) );
  FD1 data_xfi_reg_55_ ( .D(U162_Z_55), .CP(pma_tx_clk), .Q(U162_DATA3_55) );
  FD1 data_xfi_reg_56_ ( .D(U162_Z_56), .CP(pma_tx_clk), .Q(U162_DATA3_56) );
  FD1 data_xfi_reg_57_ ( .D(U162_Z_57), .CP(pma_tx_clk), .Q(U162_DATA3_57) );
  FD1 data_xfi_reg_58_ ( .D(U162_Z_58), .CP(pma_tx_clk), .Q(U162_DATA3_58) );
  FD1 data_xfi_reg_59_ ( .D(U162_Z_59), .CP(pma_tx_clk), .Q(U162_DATA3_59) );
  FD1 data_xfi_reg_60_ ( .D(U162_Z_60), .CP(pma_tx_clk), .Q(U162_DATA3_60) );
  FD1 data_xfi_reg_61_ ( .D(U162_Z_61), .CP(pma_tx_clk), .Q(U162_DATA3_61) );
  FD1 data_xfi_reg_62_ ( .D(U162_Z_62), .CP(pma_tx_clk), .Q(U162_DATA3_62) );
  FD1 data_xfi_reg_63_ ( .D(U162_Z_63), .CP(pma_tx_clk), .Q(U162_DATA3_63) );
  FD1 tx_fifo_pop_2_reg ( .D(tx_fifo_pop_pre), .CP(pma_tx_clk), .Q(
        tx_fifo_pop_2) );
  FD1 t_type_prev_reg_3_ ( .D(U160_Z_3), .CP(pma_tx_clk), .Q(n[3181]) );
  FD1 t_type_prev_reg_2_ ( .D(U160_Z_2), .CP(pma_tx_clk), .Q(n[3182]) );
  FD1 t_type_prev_reg_1_ ( .D(U160_Z_1), .CP(pma_tx_clk), .Q(n[3183]) );
  FD1 t_type_prev_reg_0_ ( .D(U160_Z_0), .CP(pma_tx_clk), .Q(n[3184]) );
  FD1 t_type_li_reg ( .D(n4900), .CP(pma_tx_clk), .Q(t_type_li) );
  FD1 tx_state_reg_3_ ( .D(U119_Z_3), .CP(pma_tx_clk), .Q(U150_DATA3_0) );
  FD1 tx_state_reg_0_ ( .D(U119_Z_0), .CP(pma_tx_clk), .Q(U153_DATA2_0) );
  FD1 tx_state_reg_2_ ( .D(U119_Z_2), .CP(pma_tx_clk), .Q(U151_DATA3_0) );
  FD1 tx_state_reg_1_ ( .D(U119_Z_1), .CP(pma_tx_clk), .Q(U152_DATA3_0) );
  FD1 tx_coded_reg_1_ ( .D(U118_Z_1), .CP(pma_tx_clk), .Q(U148_DATA3_0) );
  FD1 tx_coded_reg_0_ ( .D(U118_Z_0), .CP(pma_tx_clk), .Q(U149_DATA2_0) );
  FD1 drs1_reg ( .D(data_pat_sel), .CP(pma_tx_clk), .Q(n44) );
  FD1 drs2_reg ( .D(n44), .CP(pma_tx_clk), .Q(n97) );
  FD1 drs1_reg1 ( .D(n4399), .CP(pma_tx_clk), .Q(n41) );
  FD1 drs2_reg1 ( .D(n41), .CP(pma_tx_clk), .Q(n98) );
  FD1 test_counter_reg_0_ ( .D(U34_Z_0), .CP(pma_tx_clk), .Q(U4_DATA1_0) );
  FD1 test_counter_reg_1_ ( .D(U34_Z_1), .CP(pma_tx_clk), .Q(U4_DATA1_1) );
  FD1 test_counter_reg_2_ ( .D(U34_Z_2), .CP(pma_tx_clk), .Q(U4_DATA1_2) );
  FD1 test_counter_reg_3_ ( .D(U34_Z_3), .CP(pma_tx_clk), .Q(U4_DATA1_3) );
  FD1 test_counter_reg_4_ ( .D(U34_Z_4), .CP(pma_tx_clk), .Q(U4_DATA1_4) );
  FD1 test_counter_reg_5_ ( .D(U34_Z_5), .CP(pma_tx_clk), .Q(U4_DATA1_5) );
  FD1 test_counter_reg_6_ ( .D(U34_Z_6), .CP(pma_tx_clk), .Q(U4_DATA1_6) );
  FD1 test_counter_reg_7_ ( .D(U34_Z_7), .CP(pma_tx_clk), .Q(U4_DATA1_7) );
  FD1 test_counter_reg_8_ ( .D(U34_Z_8), .CP(pma_tx_clk), .Q(U4_DATA1_8) );
  FD1 drs1_reg2 ( .D(tx_prbs_pat_en), .CP(pma_tx_clk), .Q(n38) );
  FD1 drs2_reg2 ( .D(n38), .CP(pma_tx_clk), .Q(n4614) );
  FD1 drs1_reg3 ( .D(n4397), .CP(pma_tx_clk), .Q(n35) );
  FD1 drs2_reg3 ( .D(n35), .CP(pma_tx_clk), .Q(n4480) );
  FD1 drs1_reg4 ( .D(scr_bypass_enable), .CP(pma_tx_clk), .Q(n32) );
  FD1 drs2_reg4 ( .D(n32), .CP(pma_tx_clk), .Q(n4475) );
  FD1 tx_ts_timer_reg_8_ ( .D(U8_Z_8), .CP(pma_tx_clk), .Q(U3_U1_DATA3_8) );
  FD1 tx_ts_timer_reg_9_ ( .D(U8_Z_9), .CP(pma_tx_clk), .Q(U3_U1_DATA3_9) );
  FD1 tx_ts_timer_reg_10_ ( .D(U8_Z_10), .CP(pma_tx_clk), .Q(U3_U1_DATA3_10)
         );
  FD1 tx_ts_timer_reg_7_ ( .D(U8_Z_7), .CP(pma_tx_clk), .Q(U3_U1_DATA3_7) );
  FD1 tx_ts_timer_reg_6_ ( .D(U8_Z_6), .CP(pma_tx_clk), .Q(U3_U1_DATA3_6) );
  FD1 tx_ts_timer_reg_5_ ( .D(U8_Z_5), .CP(pma_tx_clk), .Q(U3_U1_DATA3_5) );
  FD1 tx_ts_timer_reg_4_ ( .D(U8_Z_4), .CP(pma_tx_clk), .Q(U3_U1_DATA3_4) );
  FD1 tx_ts_timer_reg_3_ ( .D(U8_Z_3), .CP(pma_tx_clk), .Q(U3_U1_DATA3_3) );
  FD1 tx_ts_timer_reg_2_ ( .D(U8_Z_2), .CP(pma_tx_clk), .Q(U3_U1_DATA3_2) );
  FD1 tx_ts_timer_reg_1_ ( .D(U8_Z_1), .CP(pma_tx_clk), .Q(U3_U1_DATA3_1) );
  FD1 tx_ts_timer_reg_0_ ( .D(U8_Z_0), .CP(pma_tx_clk), .Q(U3_U1_DATA3_0) );
  FD1 tx_lpi_state_reg_2_ ( .D(U67_Z_2), .CP(pma_tx_clk), .Q(U112_DATA3_0) );
  FD1 tx_lpi_state_reg_0_ ( .D(U67_Z_0), .CP(pma_tx_clk), .Q(U114_DATA2_0) );
  FD1 tx_lpi_state_reg_1_ ( .D(U67_Z_1), .CP(pma_tx_clk), .Q(U113_DATA3_0) );
  FD1 tx_tq_timer_reg_8_ ( .D(U7_Z_8), .CP(pma_tx_clk), .Q(sub_126_aco_A_8_)
         );
  FD1 tx_tq_timer_reg_10_ ( .D(U7_Z_10), .CP(pma_tx_clk), .Q(sub_126_aco_A_10_) );
  FD1 tx_tq_timer_reg_13_ ( .D(U7_Z_13), .CP(pma_tx_clk), .Q(sub_126_aco_A_13_) );
  FD1 tx_tq_timer_reg_14_ ( .D(U7_Z_14), .CP(pma_tx_clk), .Q(sub_126_aco_A_14_) );
  FD1 tx_tq_timer_reg_16_ ( .D(U7_Z_16), .CP(pma_tx_clk), .Q(sub_126_aco_A_16_) );
  FD1 tx_tq_timer_reg_17_ ( .D(U7_Z_17), .CP(pma_tx_clk), .Q(sub_126_aco_A_17_) );
  FD1 tx_tq_timer_reg_18_ ( .D(U7_Z_18), .CP(pma_tx_clk), .Q(sub_126_aco_A_18_) );
  FD1 tx_tq_timer_reg_19_ ( .D(U7_Z_19), .CP(pma_tx_clk), .Q(sub_126_aco_A_19_) );
  FD1 tx_tq_timer_reg_15_ ( .D(U7_Z_15), .CP(pma_tx_clk), .Q(sub_126_aco_A_15_) );
  FD1 tx_tq_timer_reg_12_ ( .D(U7_Z_12), .CP(pma_tx_clk), .Q(sub_126_aco_A_12_) );
  FD1 tx_tq_timer_reg_11_ ( .D(U7_Z_11), .CP(pma_tx_clk), .Q(sub_126_aco_A_11_) );
  FD1 tx_tq_timer_reg_9_ ( .D(U7_Z_9), .CP(pma_tx_clk), .Q(sub_126_aco_A_9_)
         );
  FD1 tx_tq_timer_reg_7_ ( .D(U7_Z_7), .CP(pma_tx_clk), .Q(sub_126_aco_A_7_)
         );
  FD1 tx_tq_timer_reg_6_ ( .D(U7_Z_6), .CP(pma_tx_clk), .Q(sub_126_aco_A_6_)
         );
  FD1 tx_tq_timer_reg_5_ ( .D(U7_Z_5), .CP(pma_tx_clk), .Q(sub_126_aco_A_5_)
         );
  FD1 tx_tq_timer_reg_4_ ( .D(U7_Z_4), .CP(pma_tx_clk), .Q(sub_126_aco_A_4_)
         );
  FD1 tx_tq_timer_reg_3_ ( .D(U7_Z_3), .CP(pma_tx_clk), .Q(sub_126_aco_A_3_)
         );
  FD1 tx_tq_timer_reg_2_ ( .D(U7_Z_2), .CP(pma_tx_clk), .Q(sub_126_aco_A_2_)
         );
  FD1 tx_tq_timer_reg_1_ ( .D(U7_Z_1), .CP(pma_tx_clk), .Q(sub_126_aco_A_1_)
         );
  FD1 tx_tq_timer_reg_0_ ( .D(U7_Z_0), .CP(pma_tx_clk), .Q(sub_126_aco_A_0_)
         );
  FD1 tx_lpi_state_reg_3_ ( .D(U67_Z_3), .CP(pma_tx_clk), .Q(U111_DATA3_0) );
  FD1 tx_refresh_timer_reg_8_ ( .D(U117_Z_8), .CP(pma_tx_clk), .Q(
        U3_U1_DATA1_8) );
  FD1 tx_refresh_timer_reg_9_ ( .D(U117_Z_9), .CP(pma_tx_clk), .Q(
        U3_U1_DATA1_9) );
  FD1 tx_refresh_timer_reg_12_ ( .D(U117_Z_12), .CP(pma_tx_clk), .Q(
        U3_U1_DATA1_12) );
  FD1 tx_refresh_timer_reg_14_ ( .D(U117_Z_14), .CP(pma_tx_clk), .Q(
        U3_U1_DATA1_14) );
  FD1 tx_refresh_timer_reg_15_ ( .D(U117_Z_15), .CP(pma_tx_clk), .Q(
        U3_U1_DATA1_15) );
  FD1 tx_refresh_timer_reg_0_ ( .D(U117_Z_0), .CP(pma_tx_clk), .Q(
        U3_U1_DATA1_0) );
  FD1 tx_refresh_timer_reg_13_ ( .D(U117_Z_13), .CP(pma_tx_clk), .Q(
        U3_U1_DATA1_13) );
  FD1 tx_refresh_timer_reg_11_ ( .D(U117_Z_11), .CP(pma_tx_clk), .Q(
        U3_U1_DATA1_11) );
  FD1 tx_refresh_timer_reg_10_ ( .D(U117_Z_10), .CP(pma_tx_clk), .Q(
        U3_U1_DATA1_10) );
  FD1 tx_refresh_timer_reg_1_ ( .D(U117_Z_1), .CP(pma_tx_clk), .Q(
        U3_U1_DATA1_1) );
  FD1 tx_refresh_timer_reg_2_ ( .D(U117_Z_2), .CP(pma_tx_clk), .Q(
        U3_U1_DATA1_2) );
  FD1 tx_refresh_timer_reg_3_ ( .D(U117_Z_3), .CP(pma_tx_clk), .Q(
        U3_U1_DATA1_3) );
  FD1 tx_refresh_timer_reg_4_ ( .D(U117_Z_4), .CP(pma_tx_clk), .Q(
        U3_U1_DATA1_4) );
  FD1 tx_refresh_timer_reg_5_ ( .D(U117_Z_5), .CP(pma_tx_clk), .Q(
        U3_U1_DATA1_5) );
  FD1 tx_refresh_timer_reg_6_ ( .D(U117_Z_6), .CP(pma_tx_clk), .Q(
        U3_U1_DATA1_6) );
  FD1 tx_refresh_timer_reg_7_ ( .D(U117_Z_7), .CP(pma_tx_clk), .Q(
        U3_U1_DATA1_7) );
  FD1 one_us_timer_reg_6_ ( .D(U5_Z_6), .CP(pma_tx_clk), .Q(sub_128_aco_A_6_)
         );
  FD1 one_us_timer_reg_7_ ( .D(U5_Z_7), .CP(pma_tx_clk), .Q(sub_128_aco_A_7_)
         );
  FD1 one_us_timer_reg_8_ ( .D(U5_Z_8), .CP(pma_tx_clk), .Q(sub_128_aco_A_8_)
         );
  FD1 tx_tw_timer_reg_8_ ( .D(U6_Z_8), .CP(pma_tx_clk), .Q(sub_127_aco_A_8_)
         );
  FD1 tx_tw_timer_reg_10_ ( .D(U6_Z_10), .CP(pma_tx_clk), .Q(sub_127_aco_A_10_) );
  FD1 tx_tw_timer_reg_11_ ( .D(U6_Z_11), .CP(pma_tx_clk), .Q(sub_127_aco_A_11_) );
  FD1 tx_tw_timer_reg_9_ ( .D(U6_Z_9), .CP(pma_tx_clk), .Q(sub_127_aco_A_9_)
         );
  FD1 tx_tw_timer_reg_0_ ( .D(U6_Z_0), .CP(pma_tx_clk), .Q(sub_127_aco_A_0_)
         );
  FD1 tx_tw_timer_reg_1_ ( .D(U6_Z_1), .CP(pma_tx_clk), .Q(sub_127_aco_A_1_)
         );
  FD1 tx_tw_timer_reg_7_ ( .D(U6_Z_7), .CP(pma_tx_clk), .Q(sub_127_aco_A_7_)
         );
  FD1 tx_tw_timer_reg_6_ ( .D(U6_Z_6), .CP(pma_tx_clk), .Q(sub_127_aco_A_6_)
         );
  FD1 tx_tw_timer_reg_5_ ( .D(U6_Z_5), .CP(pma_tx_clk), .Q(sub_127_aco_A_5_)
         );
  FD1 tx_tw_timer_reg_4_ ( .D(U6_Z_4), .CP(pma_tx_clk), .Q(sub_127_aco_A_4_)
         );
  FD1 tx_tw_timer_reg_3_ ( .D(U6_Z_3), .CP(pma_tx_clk), .Q(sub_127_aco_A_3_)
         );
  FD1 tx_tw_timer_reg_2_ ( .D(U6_Z_2), .CP(pma_tx_clk), .Q(sub_127_aco_A_2_)
         );
  FD1 one_us_timer_reg_1_ ( .D(U5_Z_1), .CP(pma_tx_clk), .Q(sub_128_aco_A_1_)
         );
  FD1 one_us_timer_reg_2_ ( .D(U5_Z_2), .CP(pma_tx_clk), .Q(sub_128_aco_A_2_)
         );
  FD1 one_us_timer_reg_3_ ( .D(U5_Z_3), .CP(pma_tx_clk), .Q(sub_128_aco_A_3_)
         );
  FD1 one_us_timer_reg_4_ ( .D(U5_Z_4), .CP(pma_tx_clk), .Q(sub_128_aco_A_4_)
         );
  FD1 one_us_timer_reg_5_ ( .D(U5_Z_5), .CP(pma_tx_clk), .Q(sub_128_aco_A_5_)
         );
  FD1 one_us_timer_reg_0_ ( .D(U5_Z_0), .CP(pma_tx_clk), .Q(sub_128_aco_A_0_)
         );
  FD1 tx_mode_reg_1_ ( .D(U66_Z_1), .CP(pma_tx_clk), .Q(tx_mode[1]) );
  FD1 tx_mode_reg_0_ ( .D(U66_Z_0), .CP(pma_tx_clk), .Q(tx_mode[0]) );
  FD1 data_prev_reg_53_ ( .D(U35_Z_53), .CP(pma_tx_clk), .Q(U37_DATA1_53) );
  FD1 data_prev_reg_47_ ( .D(U35_Z_47), .CP(pma_tx_clk), .Q(U37_DATA1_47) );
  FD1 data_prev_reg_41_ ( .D(U35_Z_41), .CP(pma_tx_clk), .Q(U37_DATA1_41) );
  FD1 data_prev_reg_35_ ( .D(U35_Z_35), .CP(pma_tx_clk), .Q(U37_DATA1_35) );
  FD1 data_prev_reg_29_ ( .D(U35_Z_29), .CP(pma_tx_clk), .Q(U37_DATA1_29) );
  FD1 data_prev_reg_23_ ( .D(U35_Z_23), .CP(pma_tx_clk), .Q(U37_DATA1_23) );
  FD1 data_prev_reg_56_ ( .D(U35_Z_56), .CP(pma_tx_clk), .Q(U37_DATA1_56) );
  FD1 data_prev_reg_50_ ( .D(U35_Z_50), .CP(pma_tx_clk), .Q(U37_DATA1_50) );
  FD1 data_prev_reg_44_ ( .D(U35_Z_44), .CP(pma_tx_clk), .Q(U37_DATA1_44) );
  FD1 data_prev_reg_19_ ( .D(U35_Z_19), .CP(pma_tx_clk), .Q(U37_DATA1_19) );
  FD1 data_prev_reg_13_ ( .D(U35_Z_13), .CP(pma_tx_clk), .Q(U37_DATA1_13) );
  FD1 data_prev_reg_7_ ( .D(U35_Z_7), .CP(pma_tx_clk), .Q(U37_DATA1_7) );
  FD1 data_prev_reg_1_ ( .D(U35_Z_1), .CP(pma_tx_clk), .Q(U37_DATA1_1) );
  FD1 data_prev_reg_40_ ( .D(U35_Z_40), .CP(pma_tx_clk), .Q(U37_DATA1_40) );
  FD1 data_prev_reg_34_ ( .D(U35_Z_34), .CP(pma_tx_clk), .Q(U37_DATA1_34) );
  FD1 data_prev_reg_28_ ( .D(U35_Z_28), .CP(pma_tx_clk), .Q(U37_DATA1_28) );
  FD1 data_prev_reg_22_ ( .D(U35_Z_22), .CP(pma_tx_clk), .Q(U37_DATA1_22) );
  FD1 data_prev_reg_16_ ( .D(U35_Z_16), .CP(pma_tx_clk), .Q(U37_DATA1_16) );
  FD1 data_prev_reg_10_ ( .D(U35_Z_10), .CP(pma_tx_clk), .Q(U37_DATA1_10) );
  FD1 data_prev_reg_4_ ( .D(U35_Z_4), .CP(pma_tx_clk), .Q(U37_DATA1_4) );
  FD1 data_prev_reg_55_ ( .D(U35_Z_55), .CP(pma_tx_clk), .Q(U37_DATA1_55) );
  FD1 data_prev_reg_49_ ( .D(U35_Z_49), .CP(pma_tx_clk), .Q(U37_DATA1_49) );
  FD1 data_prev_reg_43_ ( .D(U35_Z_43), .CP(pma_tx_clk), .Q(U37_DATA1_43) );
  FD1 data_prev_reg_37_ ( .D(U35_Z_37), .CP(pma_tx_clk), .Q(U37_DATA1_37) );
  FD1 data_prev_reg_31_ ( .D(U35_Z_31), .CP(pma_tx_clk), .Q(U37_DATA1_31) );
  FD1 data_prev_reg_25_ ( .D(U35_Z_25), .CP(pma_tx_clk), .Q(U37_DATA1_25) );
  FD1 data_prev_reg_0_ ( .D(U35_Z_0), .CP(pma_tx_clk), .Q(U37_DATA1_0) );
  FD1 data_prev_reg_52_ ( .D(U35_Z_52), .CP(pma_tx_clk), .Q(U37_DATA1_52) );
  FD1 data_prev_reg_46_ ( .D(U35_Z_46), .CP(pma_tx_clk), .Q(U37_DATA1_46) );
  FD1 data_prev_reg_39_ ( .D(U35_Z_39), .CP(pma_tx_clk), .Q(U37_DATA1_39) );
  FD1 data_prev_reg_33_ ( .D(U35_Z_33), .CP(pma_tx_clk), .Q(U37_DATA1_33) );
  FD1 data_prev_reg_27_ ( .D(U35_Z_27), .CP(pma_tx_clk), .Q(U37_DATA1_27) );
  FD1 data_prev_reg_21_ ( .D(U35_Z_21), .CP(pma_tx_clk), .Q(U37_DATA1_21) );
  FD1 data_prev_reg_15_ ( .D(U35_Z_15), .CP(pma_tx_clk), .Q(U37_DATA1_15) );
  FD1 data_prev_reg_9_ ( .D(U35_Z_9), .CP(pma_tx_clk), .Q(U37_DATA1_9) );
  FD1 data_prev_reg_3_ ( .D(U35_Z_3), .CP(pma_tx_clk), .Q(U37_DATA1_3) );
  FD1 data_prev_reg_54_ ( .D(U35_Z_54), .CP(pma_tx_clk), .Q(U37_DATA1_54) );
  FD1 data_prev_reg_48_ ( .D(U35_Z_48), .CP(pma_tx_clk), .Q(U37_DATA1_48) );
  FD1 data_prev_reg_42_ ( .D(U35_Z_42), .CP(pma_tx_clk), .Q(U37_DATA1_42) );
  FD1 data_prev_reg_17_ ( .D(U35_Z_17), .CP(pma_tx_clk), .Q(U37_DATA1_17) );
  FD1 data_prev_reg_36_ ( .D(U35_Z_36), .CP(pma_tx_clk), .Q(U37_DATA1_36) );
  FD1 data_prev_reg_11_ ( .D(U35_Z_11), .CP(pma_tx_clk), .Q(U37_DATA1_11) );
  FD1 data_prev_reg_30_ ( .D(U35_Z_30), .CP(pma_tx_clk), .Q(U37_DATA1_30) );
  FD1 data_prev_reg_5_ ( .D(U35_Z_5), .CP(pma_tx_clk), .Q(U37_DATA1_5) );
  FD1 data_prev_reg_24_ ( .D(U35_Z_24), .CP(pma_tx_clk), .Q(U37_DATA1_24) );
  FD1 data_prev_reg_18_ ( .D(U35_Z_18), .CP(pma_tx_clk), .Q(U37_DATA1_18) );
  FD1 data_prev_reg_12_ ( .D(U35_Z_12), .CP(pma_tx_clk), .Q(U37_DATA1_12) );
  FD1 data_prev_reg_6_ ( .D(U35_Z_6), .CP(pma_tx_clk), .Q(U37_DATA1_6) );
  FD1 data_prev_reg_38_ ( .D(U35_Z_38), .CP(pma_tx_clk), .Q(U37_DATA1_38) );
  FD1 data_prev_reg_57_ ( .D(U35_Z_57), .CP(pma_tx_clk), .Q(U37_DATA1_57) );
  FD1 data_prev_reg_32_ ( .D(U35_Z_32), .CP(pma_tx_clk), .Q(U37_DATA1_32) );
  FD1 data_prev_reg_51_ ( .D(U35_Z_51), .CP(pma_tx_clk), .Q(U37_DATA1_51) );
  FD1 data_prev_reg_45_ ( .D(U35_Z_45), .CP(pma_tx_clk), .Q(U37_DATA1_45) );
  FD1 data_prev_reg_26_ ( .D(U35_Z_26), .CP(pma_tx_clk), .Q(U37_DATA1_26) );
  FD1 data_prev_reg_20_ ( .D(U35_Z_20), .CP(pma_tx_clk), .Q(U37_DATA1_20) );
  FD1 data_prev_reg_14_ ( .D(U35_Z_14), .CP(pma_tx_clk), .Q(U37_DATA1_14) );
  FD1 data_prev_reg_8_ ( .D(U35_Z_8), .CP(pma_tx_clk), .Q(U37_DATA1_8) );
  FD1 data_prev_reg_2_ ( .D(U35_Z_2), .CP(pma_tx_clk), .Q(U37_DATA1_2) );
  FD1 TXxQUIET_reg ( .D(U63_Z_0), .CP(pma_tx_clk), .Q(TXxQUIET) );
  FD1 scrambler_bypass_reg ( .D(U65_Z_0), .CP(pma_tx_clk), .Q(U107_DATA1_0) );
  FD1 TXxREFRESH_reg ( .D(U64_Z_0), .CP(pma_tx_clk), .Q(TXxREFRESH) );
  IV U216 ( .A(reset_to_pma_tx), .Z(n5106) );
  IV U378 ( .A(tx_fifo_pop_pre), .Z(n5268) );
  OR2 U3546 ( .A(reset_to_pma_tx), .B(n8180), .Z(n8179) );
  AN2 U3547 ( .A(txd_xfi[9]), .B(U161_CONTROL2), .Z(n8180) );
  OR2 U3550 ( .A(reset_to_pma_tx), .B(n8183), .Z(n8182) );
  AN2 U3551 ( .A(txd_xfi[8]), .B(U161_CONTROL2), .Z(n8183) );
  AN2 U3555 ( .A(txd_xfi[7]), .B(U161_CONTROL2), .Z(n8184) );
  AN2 U3558 ( .A(txd_xfi[63]), .B(U161_CONTROL2), .Z(n8186) );
  AN2 U3561 ( .A(txd_xfi[62]), .B(U161_CONTROL2), .Z(n8188) );
  AN2 U3564 ( .A(txd_xfi[61]), .B(U161_CONTROL2), .Z(n8190) );
  AN2 U3567 ( .A(txd_xfi[60]), .B(U161_CONTROL2), .Z(n8192) );
  AN2 U3570 ( .A(txd_xfi[6]), .B(U161_CONTROL2), .Z(n8194) );
  AN2 U3573 ( .A(txd_xfi[59]), .B(U161_CONTROL2), .Z(n8196) );
  OR2 U3575 ( .A(reset_to_pma_tx), .B(n8200), .Z(n8199) );
  AN2 U3576 ( .A(txd_xfi[58]), .B(U161_CONTROL2), .Z(n8200) );
  OR2 U3579 ( .A(reset_to_pma_tx), .B(n8203), .Z(n8202) );
  AN2 U3580 ( .A(txd_xfi[57]), .B(U161_CONTROL2), .Z(n8203) );
  OR2 U3583 ( .A(reset_to_pma_tx), .B(n8206), .Z(n8205) );
  AN2 U3584 ( .A(txd_xfi[56]), .B(U161_CONTROL2), .Z(n8206) );
  AN2 U3588 ( .A(txd_xfi[55]), .B(U161_CONTROL2), .Z(n8207) );
  AN2 U3591 ( .A(txd_xfi[54]), .B(U161_CONTROL2), .Z(n8209) );
  AN2 U3594 ( .A(txd_xfi[53]), .B(U161_CONTROL2), .Z(n8211) );
  AN2 U3597 ( .A(txd_xfi[52]), .B(U161_CONTROL2), .Z(n8213) );
  AN2 U3600 ( .A(txd_xfi[51]), .B(U161_CONTROL2), .Z(n8215) );
  OR2 U3602 ( .A(reset_to_pma_tx), .B(n8219), .Z(n8218) );
  AN2 U3603 ( .A(txd_xfi[50]), .B(U161_CONTROL2), .Z(n8219) );
  AN2 U3607 ( .A(txd_xfi[5]), .B(U161_CONTROL2), .Z(n8220) );
  OR2 U3609 ( .A(reset_to_pma_tx), .B(n8224), .Z(n8223) );
  AN2 U3610 ( .A(txd_xfi[49]), .B(U161_CONTROL2), .Z(n8224) );
  OR2 U3613 ( .A(reset_to_pma_tx), .B(n8227), .Z(n8226) );
  AN2 U3614 ( .A(txd_xfi[48]), .B(U161_CONTROL2), .Z(n8227) );
  AN2 U3618 ( .A(txd_xfi[47]), .B(U161_CONTROL2), .Z(n8228) );
  AN2 U3621 ( .A(txd_xfi[46]), .B(U161_CONTROL2), .Z(n8230) );
  AN2 U3624 ( .A(txd_xfi[45]), .B(U161_CONTROL2), .Z(n8232) );
  AN2 U3627 ( .A(txd_xfi[44]), .B(U161_CONTROL2), .Z(n8234) );
  AN2 U3630 ( .A(txd_xfi[43]), .B(U161_CONTROL2), .Z(n8236) );
  OR2 U3632 ( .A(reset_to_pma_tx), .B(n8240), .Z(n8239) );
  AN2 U3633 ( .A(txd_xfi[42]), .B(U161_CONTROL2), .Z(n8240) );
  OR2 U3636 ( .A(reset_to_pma_tx), .B(n8243), .Z(n8242) );
  AN2 U3637 ( .A(txd_xfi[41]), .B(U161_CONTROL2), .Z(n8243) );
  OR2 U3640 ( .A(reset_to_pma_tx), .B(n8246), .Z(n8245) );
  AN2 U3641 ( .A(txd_xfi[40]), .B(U161_CONTROL2), .Z(n8246) );
  AN2 U3645 ( .A(txd_xfi[4]), .B(U161_CONTROL2), .Z(n8247) );
  AN2 U3648 ( .A(txd_xfi[39]), .B(U161_CONTROL2), .Z(n8249) );
  AN2 U3651 ( .A(txd_xfi[38]), .B(U161_CONTROL2), .Z(n8251) );
  AN2 U3654 ( .A(txd_xfi[37]), .B(U161_CONTROL2), .Z(n8253) );
  AN2 U3657 ( .A(txd_xfi[36]), .B(U161_CONTROL2), .Z(n8255) );
  AN2 U3660 ( .A(txd_xfi[35]), .B(U161_CONTROL2), .Z(n8257) );
  OR2 U3662 ( .A(reset_to_pma_tx), .B(n8261), .Z(n8260) );
  AN2 U3663 ( .A(txd_xfi[34]), .B(U161_CONTROL2), .Z(n8261) );
  OR2 U3666 ( .A(reset_to_pma_tx), .B(n8264), .Z(n8263) );
  AN2 U3667 ( .A(txd_xfi[33]), .B(U161_CONTROL2), .Z(n8264) );
  OR2 U3670 ( .A(reset_to_pma_tx), .B(n8267), .Z(n8266) );
  AN2 U3671 ( .A(txd_xfi[32]), .B(U161_CONTROL2), .Z(n8267) );
  AN2 U3675 ( .A(txd_xfi[31]), .B(U161_CONTROL2), .Z(n8268) );
  AN2 U3678 ( .A(txd_xfi[30]), .B(U161_CONTROL2), .Z(n8270) );
  AN2 U3681 ( .A(txd_xfi[3]), .B(U161_CONTROL2), .Z(n8272) );
  AN2 U3684 ( .A(txd_xfi[29]), .B(U161_CONTROL2), .Z(n8274) );
  AN2 U3687 ( .A(txd_xfi[28]), .B(U161_CONTROL2), .Z(n8276) );
  AN2 U3690 ( .A(txd_xfi[27]), .B(U161_CONTROL2), .Z(n8278) );
  OR2 U3692 ( .A(reset_to_pma_tx), .B(n8282), .Z(n8281) );
  AN2 U3693 ( .A(txd_xfi[26]), .B(U161_CONTROL2), .Z(n8282) );
  OR2 U3696 ( .A(reset_to_pma_tx), .B(n8285), .Z(n8284) );
  AN2 U3697 ( .A(txd_xfi[25]), .B(U161_CONTROL2), .Z(n8285) );
  OR2 U3700 ( .A(reset_to_pma_tx), .B(n8288), .Z(n8287) );
  AN2 U3701 ( .A(txd_xfi[24]), .B(U161_CONTROL2), .Z(n8288) );
  AN2 U3705 ( .A(txd_xfi[23]), .B(U161_CONTROL2), .Z(n8289) );
  AN2 U3708 ( .A(txd_xfi[22]), .B(U161_CONTROL2), .Z(n8291) );
  AN2 U3711 ( .A(txd_xfi[21]), .B(U161_CONTROL2), .Z(n8293) );
  AN2 U3714 ( .A(txd_xfi[20]), .B(U161_CONTROL2), .Z(n8295) );
  OR2 U3716 ( .A(reset_to_pma_tx), .B(n8299), .Z(n8298) );
  AN2 U3717 ( .A(txd_xfi[2]), .B(U161_CONTROL2), .Z(n8299) );
  AN2 U3721 ( .A(txd_xfi[19]), .B(U161_CONTROL2), .Z(n8300) );
  OR2 U3723 ( .A(reset_to_pma_tx), .B(n8304), .Z(n8303) );
  AN2 U3724 ( .A(txd_xfi[18]), .B(U161_CONTROL2), .Z(n8304) );
  OR2 U3727 ( .A(reset_to_pma_tx), .B(n8307), .Z(n8306) );
  AN2 U3728 ( .A(txd_xfi[17]), .B(U161_CONTROL2), .Z(n8307) );
  OR2 U3731 ( .A(reset_to_pma_tx), .B(n8310), .Z(n8309) );
  AN2 U3732 ( .A(txd_xfi[16]), .B(U161_CONTROL2), .Z(n8310) );
  AN2 U3736 ( .A(txd_xfi[15]), .B(U161_CONTROL2), .Z(n8311) );
  AN2 U3739 ( .A(txd_xfi[14]), .B(U161_CONTROL2), .Z(n8313) );
  AN2 U3742 ( .A(txd_xfi[13]), .B(U161_CONTROL2), .Z(n8315) );
  AN2 U3745 ( .A(txd_xfi[12]), .B(U161_CONTROL2), .Z(n8317) );
  AN2 U3748 ( .A(txd_xfi[11]), .B(U161_CONTROL2), .Z(n8319) );
  OR2 U3750 ( .A(reset_to_pma_tx), .B(n8323), .Z(n8322) );
  AN2 U3751 ( .A(txd_xfi[10]), .B(U161_CONTROL2), .Z(n8323) );
  OR2 U3754 ( .A(reset_to_pma_tx), .B(n8326), .Z(n8325) );
  AN2 U3755 ( .A(txd_xfi[1]), .B(U161_CONTROL2), .Z(n8326) );
  OR2 U3758 ( .A(reset_to_pma_tx), .B(n8329), .Z(n8328) );
  AN2 U3759 ( .A(txd_xfi[0]), .B(U161_CONTROL2), .Z(n8329) );
  OR2 U3762 ( .A(reset_to_pma_tx), .B(n8332), .Z(n8331) );
  AN2 U3763 ( .A(txc_xfi[7]), .B(U161_CONTROL2), .Z(n8332) );
  OR2 U3766 ( .A(reset_to_pma_tx), .B(n8335), .Z(n8334) );
  AN2 U3767 ( .A(txc_xfi[6]), .B(U161_CONTROL2), .Z(n8335) );
  OR2 U3770 ( .A(reset_to_pma_tx), .B(n8338), .Z(n8337) );
  AN2 U3771 ( .A(txc_xfi[5]), .B(U161_CONTROL2), .Z(n8338) );
  OR2 U3774 ( .A(reset_to_pma_tx), .B(n8341), .Z(n8340) );
  AN2 U3775 ( .A(txc_xfi[4]), .B(U161_CONTROL2), .Z(n8341) );
  OR2 U3778 ( .A(reset_to_pma_tx), .B(n8344), .Z(n8343) );
  AN2 U3779 ( .A(txc_xfi[3]), .B(U161_CONTROL2), .Z(n8344) );
  OR2 U3782 ( .A(reset_to_pma_tx), .B(n8347), .Z(n8346) );
  AN2 U3783 ( .A(txc_xfi[2]), .B(U161_CONTROL2), .Z(n8347) );
  OR2 U3786 ( .A(reset_to_pma_tx), .B(n8350), .Z(n8349) );
  AN2 U3787 ( .A(txc_xfi[1]), .B(U161_CONTROL2), .Z(n8350) );
  OR2 U3790 ( .A(reset_to_pma_tx), .B(n8353), .Z(n8352) );
  AN2 U3791 ( .A(txc_xfi[0]), .B(U161_CONTROL2), .Z(n8353) );
  AN2 U3793 ( .A(n5268), .B(n5106), .Z(U161_CONTROL3) );
  AN2 U3794 ( .A(n5106), .B(tx_fifo_pop_pre), .Z(U161_CONTROL2) );
  AN2 U4189 ( .A(n8647), .B(n1235), .Z(n940) );
  AN2 U4190 ( .A(n1226), .B(n8648), .Z(n8647) );
  IV U4191 ( .A(n5270), .Z(n8642) );
  IV U4192 ( .A(n5261), .Z(n8641) );
  AN2 U4193 ( .A(n8649), .B(n8650), .Z(n817) );
  AN2 U4194 ( .A(n5627), .B(n8651), .Z(n8649) );
  AN2 U4195 ( .A(n97), .B(n8650), .Z(n816) );
  AN2 U4196 ( .A(n8652), .B(n8650), .Z(n750) );
  IV U4197 ( .A(n8653), .Z(n8650) );
  OR2 U4198 ( .A(n749), .B(n5684), .Z(n8653) );
  AN2 U4199 ( .A(U4_DATA1_7), .B(n8651), .Z(n8652) );
  IV U4200 ( .A(n97), .Z(n8651) );
  IV U4201 ( .A(n4475), .Z(n5685) );
  IV U4202 ( .A(U111_DATA3_0), .Z(n5527) );
  IV U4203 ( .A(U112_DATA3_0), .Z(n5526) );
  IV U4204 ( .A(U113_DATA3_0), .Z(n5525) );
  IV U4205 ( .A(n8654), .Z(n5521) );
  OR2 U4206 ( .A(n2576), .B(n2575), .Z(n8654) );
  IV U4207 ( .A(n8655), .Z(n5520) );
  OR2 U4208 ( .A(n2579), .B(n2578), .Z(n8655) );
  IV U4209 ( .A(n8656), .Z(n5519) );
  OR2 U4210 ( .A(n2582), .B(n2581), .Z(n8656) );
  IV U4211 ( .A(n8657), .Z(n5518) );
  OR2 U4212 ( .A(n2585), .B(n2584), .Z(n8657) );
  IV U4213 ( .A(U114_DATA2_0), .Z(n5517) );
  IV U4214 ( .A(n8658), .Z(n5515) );
  OR2 U4215 ( .A(n8659), .B(n8660), .Z(n8658) );
  AN2 U4216 ( .A(n8661), .B(U3_U1_DATA1_0), .Z(n8660) );
  AN2 U4217 ( .A(n8662), .B(U3_U1_DATA3_0), .Z(n8659) );
  IV U4218 ( .A(r224_GTV2_1_), .Z(n5514) );
  IV U4219 ( .A(r224_GTV_2_), .Z(n5513) );
  IV U4220 ( .A(r224_GTV2_2_), .Z(n5512) );
  IV U4221 ( .A(r224_GTV_3_), .Z(n5511) );
  IV U4222 ( .A(r224_GTV2_3_), .Z(n5510) );
  IV U4223 ( .A(r224_GTV_4_), .Z(n5509) );
  IV U4224 ( .A(r224_GTV2_4_), .Z(n5508) );
  IV U4225 ( .A(r224_GTV_5_), .Z(n5507) );
  IV U4226 ( .A(r224_GTV2_5_), .Z(n5506) );
  IV U4227 ( .A(r224_GTV_6_), .Z(n5505) );
  IV U4228 ( .A(r224_GTV2_6_), .Z(n5504) );
  IV U4229 ( .A(r224_GTV_7_), .Z(n5503) );
  IV U4230 ( .A(r224_GTV2_7_), .Z(n5502) );
  IV U4231 ( .A(r224_GTV_8_), .Z(n5501) );
  IV U4232 ( .A(r224_GTV2_8_), .Z(n5500) );
  IV U4233 ( .A(r224_GTV_9_), .Z(n5499) );
  IV U4234 ( .A(r224_GTV2_9_), .Z(n5498) );
  IV U4235 ( .A(r224_GTV_10_), .Z(n5497) );
  IV U4236 ( .A(r224_GTV2_10_), .Z(n5496) );
  IV U4237 ( .A(r224_GTV_11_), .Z(n5495) );
  IV U4238 ( .A(r224_GTV2_11_), .Z(n5494) );
  IV U4239 ( .A(r224_GTV_12_), .Z(n5493) );
  IV U4240 ( .A(r224_GTV2_12_), .Z(n5492) );
  IV U4241 ( .A(r224_GTV_13_), .Z(n5491) );
  IV U4242 ( .A(r224_GTV2_13_), .Z(n5490) );
  IV U4243 ( .A(r224_GTV_14_), .Z(n5489) );
  IV U4244 ( .A(r224_GTV2_14_), .Z(n5488) );
  IV U4245 ( .A(r224_GTV_15_), .Z(n5487) );
  IV U4246 ( .A(r224_GTV2_15_), .Z(n5486) );
  IV U4247 ( .A(r224_GT), .Z(n5485) );
  IV U4248 ( .A(n8663), .Z(n5481) );
  OR2 U4249 ( .A(n2564), .B(n2563), .Z(n8663) );
  IV U4250 ( .A(n8664), .Z(n5480) );
  OR2 U4251 ( .A(n2567), .B(n2566), .Z(n8664) );
  IV U4252 ( .A(n8665), .Z(n5479) );
  OR2 U4253 ( .A(n2570), .B(n2569), .Z(n8665) );
  IV U4254 ( .A(n8666), .Z(n5478) );
  OR2 U4255 ( .A(n2573), .B(n2572), .Z(n8666) );
  IV U4256 ( .A(tx_mode[1]), .Z(n5477) );
  IV U4257 ( .A(n4369), .Z(n5476) );
  IV U4258 ( .A(tx_mode[0]), .Z(n5474) );
  IV U4259 ( .A(U150_DATA3_0), .Z(n5471) );
  IV U4260 ( .A(U151_DATA3_0), .Z(n5470) );
  IV U4261 ( .A(U152_DATA3_0), .Z(n5469) );
  IV U4262 ( .A(U153_DATA2_0), .Z(n5467) );
  IV U4263 ( .A(U148_DATA3_0), .Z(n5462) );
  IV U4264 ( .A(U149_DATA2_0), .Z(n5459) );
  IV U4265 ( .A(n[3182]), .Z(n5455) );
  IV U4266 ( .A(n[3183]), .Z(n5454) );
  IV U4267 ( .A(n3521), .Z(n5453) );
  IV U4268 ( .A(U156_Z_33), .Z(n5451) );
  IV U4269 ( .A(U156_Z_32), .Z(n5450) );
  IV U4270 ( .A(U156_Z_31), .Z(n5449) );
  IV U4271 ( .A(U156_Z_30), .Z(n5448) );
  IV U4272 ( .A(U156_Z_29), .Z(n5447) );
  IV U4273 ( .A(n8667), .Z(n5446) );
  IV U4274 ( .A(U158_Z_14), .Z(n5445) );
  IV U4275 ( .A(U158_Z_13), .Z(n5437) );
  IV U4276 ( .A(n1806), .Z(n5435) );
  IV U4277 ( .A(n1825), .Z(n5434) );
  IV U4278 ( .A(U156_Z_28), .Z(n5433) );
  IV U4279 ( .A(U156_Z_27), .Z(n5432) );
  IV U4280 ( .A(U156_Z_26), .Z(n5431) );
  IV U4281 ( .A(U156_Z_25), .Z(n5430) );
  IV U4282 ( .A(U156_Z_24), .Z(n5429) );
  IV U4283 ( .A(n8668), .Z(n5428) );
  IV U4284 ( .A(U158_Z_11), .Z(n5427) );
  IV U4285 ( .A(U159_Z_7), .Z(n5419) );
  IV U4286 ( .A(n1812), .Z(n5417) );
  IV U4287 ( .A(n1828), .Z(n5416) );
  IV U4288 ( .A(U156_Z_23), .Z(n5415) );
  IV U4289 ( .A(U156_Z_22), .Z(n5414) );
  IV U4290 ( .A(U156_Z_21), .Z(n5413) );
  IV U4291 ( .A(U156_Z_20), .Z(n5412) );
  IV U4292 ( .A(U156_Z_19), .Z(n5411) );
  IV U4293 ( .A(n8669), .Z(n5410) );
  IV U4294 ( .A(U158_Z_9), .Z(n5409) );
  IV U4295 ( .A(U159_Z_6), .Z(n5401) );
  IV U4296 ( .A(n1818), .Z(n5399) );
  IV U4297 ( .A(n1831), .Z(n5398) );
  IV U4298 ( .A(U157_Z_5), .Z(n5397) );
  IV U4299 ( .A(U156_Z_18), .Z(n5396) );
  IV U4300 ( .A(U156_Z_17), .Z(n5395) );
  IV U4301 ( .A(U157_Z_4), .Z(n5394) );
  IV U4302 ( .A(U157_Z_3), .Z(n5393) );
  IV U4303 ( .A(U159_Z_5), .Z(n5392) );
  IV U4304 ( .A(U158_Z_8), .Z(n5391) );
  IV U4305 ( .A(n1349), .Z(n5390) );
  IV U4306 ( .A(n1868), .Z(n5382) );
  IV U4307 ( .A(U159_Z_4), .Z(n5381) );
  IV U4308 ( .A(n1821), .Z(n5379) );
  IV U4309 ( .A(n1834), .Z(n5378) );
  IV U4310 ( .A(n1861), .Z(n5377) );
  IV U4311 ( .A(U156_Z_16), .Z(n5376) );
  IV U4312 ( .A(U156_Z_15), .Z(n5375) );
  IV U4313 ( .A(U156_Z_14), .Z(n5374) );
  IV U4314 ( .A(U156_Z_13), .Z(n5373) );
  IV U4315 ( .A(U156_Z_12), .Z(n5372) );
  IV U4316 ( .A(n8670), .Z(n5371) );
  IV U4317 ( .A(U158_Z_6), .Z(n5370) );
  IV U4318 ( .A(U158_Z_5), .Z(n5362) );
  IV U4319 ( .A(n1800), .Z(n5360) );
  IV U4320 ( .A(n1837), .Z(n5359) );
  IV U4321 ( .A(U156_Z_11), .Z(n5358) );
  IV U4322 ( .A(U156_Z_10), .Z(n5357) );
  IV U4323 ( .A(U156_Z_9), .Z(n5356) );
  IV U4324 ( .A(U156_Z_8), .Z(n5355) );
  IV U4325 ( .A(U156_Z_7), .Z(n5354) );
  IV U4326 ( .A(n8671), .Z(n5353) );
  IV U4327 ( .A(U158_Z_3), .Z(n5352) );
  IV U4328 ( .A(U159_Z_3), .Z(n5344) );
  IV U4329 ( .A(n1803), .Z(n5342) );
  IV U4330 ( .A(n1840), .Z(n5341) );
  IV U4331 ( .A(U156_Z_6), .Z(n5340) );
  IV U4332 ( .A(U156_Z_5), .Z(n5339) );
  IV U4333 ( .A(U156_Z_4), .Z(n5338) );
  IV U4334 ( .A(U156_Z_3), .Z(n5337) );
  IV U4335 ( .A(U156_Z_2), .Z(n5336) );
  IV U4336 ( .A(n8672), .Z(n5335) );
  IV U4337 ( .A(U158_Z_1), .Z(n5334) );
  IV U4338 ( .A(U159_Z_2), .Z(n5326) );
  IV U4339 ( .A(n1809), .Z(n5324) );
  IV U4340 ( .A(n1843), .Z(n5323) );
  IV U4341 ( .A(U157_Z_2), .Z(n5322) );
  IV U4342 ( .A(U156_Z_1), .Z(n5321) );
  IV U4343 ( .A(U156_Z_0), .Z(n5320) );
  IV U4344 ( .A(U157_Z_1), .Z(n5319) );
  IV U4345 ( .A(U157_Z_0), .Z(n5318) );
  IV U4346 ( .A(U159_Z_1), .Z(n5317) );
  IV U4347 ( .A(U158_Z_0), .Z(n5316) );
  IV U4348 ( .A(n1268), .Z(n5315) );
  IV U4349 ( .A(n1857), .Z(n5307) );
  IV U4350 ( .A(U159_Z_0), .Z(n5306) );
  IV U4351 ( .A(n1815), .Z(n5304) );
  IV U4352 ( .A(n1846), .Z(n5303) );
  IV U4353 ( .A(n1850), .Z(n5302) );
  IV U4354 ( .A(U154_Z_5), .Z(n5301) );
  IV U4355 ( .A(U154_Z_4), .Z(n5300) );
  IV U4356 ( .A(U154_Z_3), .Z(n5299) );
  IV U4357 ( .A(U155_Z_1), .Z(n5298) );
  IV U4358 ( .A(U154_Z_2), .Z(n5297) );
  IV U4359 ( .A(U154_Z_1), .Z(n5296) );
  IV U4360 ( .A(U154_Z_0), .Z(n5295) );
  IV U4361 ( .A(n1506), .Z(n5294) );
  IV U4362 ( .A(n8644), .Z(n5288) );
  OR2 U4363 ( .A(n126), .B(n8673), .Z(n8644) );
  IV U4364 ( .A(n336), .Z(n5285) );
  IV U4365 ( .A(n8646), .Z(n5284) );
  OR2 U4366 ( .A(n8674), .B(n8675), .Z(n8646) );
  IV U4367 ( .A(n331), .Z(n5282) );
  IV U4368 ( .A(n8643), .Z(n5281) );
  OR2 U4369 ( .A(n8676), .B(n8677), .Z(n8643) );
  IV U4370 ( .A(n314), .Z(n8677) );
  IV U4371 ( .A(n8645), .Z(n5279) );
  OR2 U4372 ( .A(n8678), .B(n8679), .Z(n8645) );
  IV U4373 ( .A(n311), .Z(n8679) );
  IV U4374 ( .A(n334), .Z(n5277) );
  IV U4375 ( .A(n4372), .Z(n5275) );
  IV U4376 ( .A(U155_Z_0), .Z(n5274) );
  AN2 U4377 ( .A(n8680), .B(n315), .Z(n5270) );
  IV U4378 ( .A(n328), .Z(n5269) );
  IV U4379 ( .A(n325), .Z(n5264) );
  IV U4380 ( .A(n324), .Z(n5263) );
  AN2 U4381 ( .A(n8681), .B(n8682), .Z(n5261) );
  AN2 U4382 ( .A(n8683), .B(n322), .Z(n8682) );
  IV U4383 ( .A(n8684), .Z(n8681) );
  OR2 U4384 ( .A(n321), .B(n320), .Z(n8684) );
  IV U4385 ( .A(n326), .Z(n5259) );
  IV U4386 ( .A(n327), .Z(n5236) );
  IV U4387 ( .A(U161_Z_0), .Z(n5105) );
  IV U4388 ( .A(U161_Z_1), .Z(n5104) );
  IV U4389 ( .A(U161_Z_2), .Z(n5103) );
  IV U4390 ( .A(n3479), .Z(n5102) );
  IV U4391 ( .A(U161_Z_3), .Z(n5101) );
  IV U4392 ( .A(U161_Z_4), .Z(n5100) );
  IV U4393 ( .A(U161_Z_5), .Z(n5099) );
  IV U4394 ( .A(U161_Z_6), .Z(n5098) );
  IV U4395 ( .A(n3419), .Z(n5097) );
  IV U4396 ( .A(n3433), .Z(n5096) );
  IV U4397 ( .A(n3499), .Z(n5095) );
  IV U4398 ( .A(U161_Z_7), .Z(n5094) );
  IV U4399 ( .A(U162_Z_0), .Z(n5093) );
  IV U4400 ( .A(U162_Z_1), .Z(n5092) );
  IV U4401 ( .A(U162_Z_10), .Z(n5091) );
  IV U4402 ( .A(U162_Z_11), .Z(n5090) );
  IV U4403 ( .A(U162_Z_12), .Z(n5089) );
  IV U4404 ( .A(U162_Z_13), .Z(n5088) );
  IV U4405 ( .A(U162_Z_14), .Z(n5087) );
  IV U4406 ( .A(U162_Z_15), .Z(n5086) );
  IV U4407 ( .A(U162_Z_16), .Z(n5085) );
  IV U4408 ( .A(U162_Z_17), .Z(n5084) );
  IV U4409 ( .A(U162_Z_18), .Z(n5083) );
  IV U4410 ( .A(U162_Z_19), .Z(n5082) );
  IV U4411 ( .A(U162_Z_2), .Z(n5081) );
  IV U4412 ( .A(U162_Z_20), .Z(n5080) );
  IV U4413 ( .A(U162_Z_21), .Z(n5079) );
  IV U4414 ( .A(U162_Z_22), .Z(n5078) );
  IV U4415 ( .A(n3547), .Z(n5077) );
  IV U4416 ( .A(n3222), .Z(n5076) );
  IV U4417 ( .A(n4031), .Z(n5075) );
  IV U4418 ( .A(n4039), .Z(n5074) );
  IV U4419 ( .A(n4047), .Z(n5073) );
  IV U4420 ( .A(n4063), .Z(n5072) );
  IV U4421 ( .A(n4087), .Z(n5071) );
  IV U4422 ( .A(U162_Z_23), .Z(n5070) );
  IV U4423 ( .A(n3335), .Z(n5069) );
  IV U4424 ( .A(n4055), .Z(n5068) );
  IV U4425 ( .A(n4071), .Z(n5067) );
  IV U4426 ( .A(n4079), .Z(n5066) );
  IV U4427 ( .A(n4095), .Z(n5065) );
  IV U4428 ( .A(U162_Z_24), .Z(n5064) );
  IV U4429 ( .A(U162_Z_25), .Z(n5063) );
  IV U4430 ( .A(U162_Z_26), .Z(n5062) );
  IV U4431 ( .A(U162_Z_27), .Z(n5061) );
  IV U4432 ( .A(U162_Z_28), .Z(n5060) );
  IV U4433 ( .A(U162_Z_29), .Z(n5059) );
  IV U4434 ( .A(U162_Z_3), .Z(n5058) );
  IV U4435 ( .A(U162_Z_30), .Z(n5057) );
  IV U4436 ( .A(n3556), .Z(n5056) );
  IV U4437 ( .A(n3221), .Z(n5055) );
  IV U4438 ( .A(n4103), .Z(n5054) );
  IV U4439 ( .A(n4111), .Z(n5053) );
  IV U4440 ( .A(n4119), .Z(n5052) );
  IV U4441 ( .A(n4135), .Z(n5051) );
  IV U4442 ( .A(n4159), .Z(n5050) );
  IV U4443 ( .A(U162_Z_31), .Z(n5049) );
  IV U4444 ( .A(n3410), .Z(n5048) );
  IV U4445 ( .A(n4127), .Z(n5047) );
  IV U4446 ( .A(n4143), .Z(n5046) );
  IV U4447 ( .A(n4151), .Z(n5045) );
  IV U4448 ( .A(n4167), .Z(n5044) );
  IV U4449 ( .A(U162_Z_32), .Z(n5043) );
  IV U4450 ( .A(U162_Z_33), .Z(n5042) );
  IV U4451 ( .A(U162_Z_34), .Z(n5041) );
  IV U4452 ( .A(U162_Z_35), .Z(n5040) );
  IV U4453 ( .A(U162_Z_36), .Z(n5039) );
  IV U4454 ( .A(U162_Z_37), .Z(n5038) );
  IV U4455 ( .A(U162_Z_38), .Z(n5037) );
  IV U4456 ( .A(n3515), .Z(n5036) );
  IV U4457 ( .A(n3564), .Z(n5035) );
  IV U4458 ( .A(n3220), .Z(n5034) );
  IV U4459 ( .A(n3599), .Z(n5033) );
  IV U4460 ( .A(n3607), .Z(n5032) );
  IV U4461 ( .A(n3615), .Z(n5031) );
  IV U4462 ( .A(n3631), .Z(n5030) );
  IV U4463 ( .A(n3655), .Z(n5029) );
  IV U4464 ( .A(U162_Z_39), .Z(n5028) );
  IV U4465 ( .A(n3350), .Z(n5027) );
  IV U4466 ( .A(n3442), .Z(n5026) );
  IV U4467 ( .A(n3507), .Z(n5025) );
  IV U4468 ( .A(n3623), .Z(n5024) );
  IV U4469 ( .A(n3639), .Z(n5023) );
  IV U4470 ( .A(n3647), .Z(n5022) );
  IV U4471 ( .A(n3663), .Z(n5021) );
  IV U4472 ( .A(U162_Z_4), .Z(n5020) );
  IV U4473 ( .A(U162_Z_40), .Z(n5019) );
  IV U4474 ( .A(U162_Z_41), .Z(n5018) );
  IV U4475 ( .A(U162_Z_42), .Z(n5017) );
  IV U4476 ( .A(U162_Z_43), .Z(n5016) );
  IV U4477 ( .A(U162_Z_44), .Z(n5015) );
  IV U4478 ( .A(U162_Z_45), .Z(n5014) );
  IV U4479 ( .A(U162_Z_46), .Z(n5013) );
  IV U4480 ( .A(n3573), .Z(n5012) );
  IV U4481 ( .A(n3219), .Z(n5011) );
  IV U4482 ( .A(n3671), .Z(n5010) );
  IV U4483 ( .A(n3679), .Z(n5009) );
  IV U4484 ( .A(n3687), .Z(n5008) );
  IV U4485 ( .A(n3703), .Z(n5007) );
  IV U4486 ( .A(n3727), .Z(n5006) );
  IV U4487 ( .A(U162_Z_47), .Z(n5005) );
  IV U4488 ( .A(n3365), .Z(n5004) );
  IV U4489 ( .A(n3695), .Z(n5003) );
  IV U4490 ( .A(n3711), .Z(n5002) );
  IV U4491 ( .A(n3719), .Z(n5001) );
  IV U4492 ( .A(n3735), .Z(n5000) );
  IV U4493 ( .A(U162_Z_48), .Z(n4999) );
  IV U4494 ( .A(U162_Z_49), .Z(n4998) );
  IV U4495 ( .A(U162_Z_5), .Z(n4997) );
  IV U4496 ( .A(U162_Z_50), .Z(n4996) );
  IV U4497 ( .A(U162_Z_51), .Z(n4995) );
  IV U4498 ( .A(U162_Z_52), .Z(n4994) );
  IV U4499 ( .A(U162_Z_53), .Z(n4993) );
  IV U4500 ( .A(U162_Z_54), .Z(n4992) );
  IV U4501 ( .A(n3582), .Z(n4991) );
  IV U4502 ( .A(n3218), .Z(n4990) );
  IV U4503 ( .A(n3743), .Z(n4989) );
  IV U4504 ( .A(n3751), .Z(n4988) );
  IV U4505 ( .A(n3759), .Z(n4987) );
  IV U4506 ( .A(n3775), .Z(n4986) );
  IV U4507 ( .A(n3799), .Z(n4985) );
  IV U4508 ( .A(U162_Z_55), .Z(n4984) );
  IV U4509 ( .A(n3380), .Z(n4983) );
  IV U4510 ( .A(n3767), .Z(n4982) );
  IV U4511 ( .A(n3783), .Z(n4981) );
  IV U4512 ( .A(n3791), .Z(n4980) );
  IV U4513 ( .A(n3807), .Z(n4979) );
  IV U4514 ( .A(U162_Z_56), .Z(n4978) );
  IV U4515 ( .A(U162_Z_57), .Z(n4977) );
  IV U4516 ( .A(U162_Z_58), .Z(n4976) );
  IV U4517 ( .A(U162_Z_59), .Z(n4975) );
  IV U4518 ( .A(U162_Z_6), .Z(n4974) );
  IV U4519 ( .A(U162_Z_60), .Z(n4973) );
  IV U4520 ( .A(U162_Z_61), .Z(n4972) );
  IV U4521 ( .A(U162_Z_62), .Z(n4971) );
  IV U4522 ( .A(n3591), .Z(n4970) );
  IV U4523 ( .A(n3217), .Z(n4969) );
  IV U4524 ( .A(n3815), .Z(n4968) );
  IV U4525 ( .A(n3823), .Z(n4967) );
  IV U4526 ( .A(n3831), .Z(n4966) );
  IV U4527 ( .A(n3847), .Z(n4965) );
  IV U4528 ( .A(n3871), .Z(n4964) );
  IV U4529 ( .A(U162_Z_63), .Z(n4963) );
  IV U4530 ( .A(n3395), .Z(n4962) );
  IV U4531 ( .A(n3839), .Z(n4961) );
  IV U4532 ( .A(n3855), .Z(n4960) );
  IV U4533 ( .A(n3863), .Z(n4959) );
  IV U4534 ( .A(n3879), .Z(n4958) );
  IV U4535 ( .A(n3495), .Z(n4957) );
  IV U4536 ( .A(n3529), .Z(n4956) );
  IV U4537 ( .A(n3224), .Z(n4955) );
  IV U4538 ( .A(n3887), .Z(n4954) );
  IV U4539 ( .A(n3895), .Z(n4953) );
  IV U4540 ( .A(n3903), .Z(n4952) );
  IV U4541 ( .A(n3919), .Z(n4951) );
  IV U4542 ( .A(n3943), .Z(n4950) );
  IV U4543 ( .A(U162_Z_7), .Z(n4949) );
  IV U4544 ( .A(n3305), .Z(n4948) );
  IV U4545 ( .A(n3428), .Z(n4947) );
  IV U4546 ( .A(n3487), .Z(n4946) );
  IV U4547 ( .A(n3911), .Z(n4945) );
  IV U4548 ( .A(n3927), .Z(n4944) );
  IV U4549 ( .A(n3935), .Z(n4943) );
  IV U4550 ( .A(n3951), .Z(n4942) );
  IV U4551 ( .A(U162_Z_8), .Z(n4941) );
  IV U4552 ( .A(n3320), .Z(n4940) );
  IV U4553 ( .A(n3967), .Z(n4939) );
  IV U4554 ( .A(n3975), .Z(n4938) );
  IV U4555 ( .A(n3983), .Z(n4937) );
  IV U4556 ( .A(n3991), .Z(n4936) );
  IV U4557 ( .A(n3999), .Z(n4935) );
  IV U4558 ( .A(U162_Z_9), .Z(n4934) );
  IV U4559 ( .A(n3538), .Z(n4933) );
  IV U4560 ( .A(n3450), .Z(n4932) );
  IV U4561 ( .A(n3462), .Z(n4931) );
  IV U4562 ( .A(n3223), .Z(n4929) );
  IV U4563 ( .A(n3474), .Z(n4928) );
  IV U4564 ( .A(n3959), .Z(n4927) );
  IV U4565 ( .A(n4007), .Z(n4926) );
  IV U4566 ( .A(n4015), .Z(n4925) );
  IV U4567 ( .A(n4023), .Z(n4924) );
  IV U4568 ( .A(U160_DATA2_1), .Z(n4918) );
  IV U4569 ( .A(U160_DATA2_0), .Z(n4917) );
  IV U4570 ( .A(U160_DATA2_2), .Z(n4913) );
  IV U4571 ( .A(n2964), .Z(n4911) );
  AN2 U4572 ( .A(n8685), .B(n318), .Z(n339) );
  AN2 U4573 ( .A(n8686), .B(n8687), .Z(n8685) );
  IV U4574 ( .A(n317), .Z(n8687) );
  AN2 U4575 ( .A(n317), .B(n8686), .Z(n338) );
  AN2 U4576 ( .A(n308), .B(n8688), .Z(n336) );
  AN2 U4577 ( .A(n8673), .B(n8689), .Z(n8688) );
  IV U4578 ( .A(n126), .Z(n8689) );
  IV U4579 ( .A(n307), .Z(n8673) );
  IV U4580 ( .A(n5276), .Z(n335) );
  OR2 U4581 ( .A(n8690), .B(n8691), .Z(n5276) );
  AN2 U4582 ( .A(n310), .B(n8692), .Z(n334) );
  AN2 U4583 ( .A(n8691), .B(n8693), .Z(n8692) );
  IV U4584 ( .A(n8690), .Z(n8693) );
  IV U4585 ( .A(n309), .Z(n8691) );
  AN2 U4586 ( .A(n313), .B(n8694), .Z(n331) );
  AN2 U4587 ( .A(n8675), .B(n8695), .Z(n8694) );
  IV U4588 ( .A(n8674), .Z(n8695) );
  IV U4589 ( .A(n312), .Z(n8675) );
  AN2 U4590 ( .A(n316), .B(n8696), .Z(n328) );
  IV U4591 ( .A(n8697), .Z(n8696) );
  OR2 U4592 ( .A(n315), .B(n8698), .Z(n8697) );
  AN2 U4593 ( .A(n8699), .B(n3290), .Z(n3268) );
  IV U4594 ( .A(n8700), .Z(n8699) );
  OR2 U4595 ( .A(n8701), .B(n3281), .Z(n8700) );
  AN2 U4596 ( .A(n3290), .B(n8701), .Z(n3267) );
  IV U4597 ( .A(n3288), .Z(n8701) );
  AN2 U4598 ( .A(n8702), .B(n319), .Z(n326) );
  AN2 U4599 ( .A(n8683), .B(n320), .Z(n325) );
  AN2 U4600 ( .A(n321), .B(n8703), .Z(n324) );
  AN2 U4601 ( .A(n8704), .B(n8683), .Z(n8703) );
  AN2 U4602 ( .A(n8705), .B(n8702), .Z(n8683) );
  AN2 U4603 ( .A(n8686), .B(n8706), .Z(n8702) );
  IV U4604 ( .A(n8707), .Z(n8706) );
  OR2 U4605 ( .A(n318), .B(n317), .Z(n8707) );
  AN2 U4606 ( .A(n8680), .B(n8708), .Z(n8686) );
  IV U4607 ( .A(n8709), .Z(n8708) );
  OR2 U4608 ( .A(n316), .B(n315), .Z(n8709) );
  IV U4609 ( .A(n8698), .Z(n8680) );
  OR2 U4610 ( .A(n314), .B(n8676), .Z(n8698) );
  OR2 U4611 ( .A(n8674), .B(n8710), .Z(n8676) );
  OR2 U4612 ( .A(n313), .B(n312), .Z(n8710) );
  OR2 U4613 ( .A(n311), .B(n8678), .Z(n8674) );
  OR2 U4614 ( .A(n8690), .B(n8711), .Z(n8678) );
  OR2 U4615 ( .A(n310), .B(n309), .Z(n8711) );
  OR2 U4616 ( .A(n126), .B(n8712), .Z(n8690) );
  OR2 U4617 ( .A(n308), .B(n307), .Z(n8712) );
  IV U4618 ( .A(n319), .Z(n8705) );
  IV U4619 ( .A(n320), .Z(n8704) );
  OR2 U4620 ( .A(n8713), .B(n8714), .Z(n2774) );
  OR2 U4621 ( .A(n8715), .B(n8716), .Z(n8714) );
  AN2 U4622 ( .A(n2534), .B(n2533), .Z(n8716) );
  OR2 U4623 ( .A(n8717), .B(n8718), .Z(n8713) );
  OR2 U4624 ( .A(n8719), .B(n8662), .Z(n8718) );
  AN2 U4625 ( .A(n8720), .B(n8721), .Z(n239) );
  AN2 U4626 ( .A(n1397), .B(n1298), .Z(n8720) );
  AN2 U4627 ( .A(n8722), .B(n8723), .Z(n223) );
  AN2 U4628 ( .A(n1423), .B(n1318), .Z(n8722) );
  AN2 U4629 ( .A(n8724), .B(n8725), .Z(n207) );
  AN2 U4630 ( .A(n1446), .B(n1337), .Z(n8724) );
  AN2 U4631 ( .A(n8726), .B(n8727), .Z(n191) );
  AN2 U4632 ( .A(n1456), .B(n1358), .Z(n8726) );
  OR2 U4633 ( .A(n8728), .B(n8729), .Z(n1909) );
  OR2 U4634 ( .A(n1929), .B(n5249), .Z(n8729) );
  OR2 U4635 ( .A(n5247), .B(n8730), .Z(n1905) );
  OR2 U4636 ( .A(n8731), .B(n8730), .Z(n1901) );
  OR2 U4637 ( .A(n8732), .B(n8733), .Z(n8730) );
  OR2 U4638 ( .A(n8734), .B(n8728), .Z(n8733) );
  OR2 U4639 ( .A(n5248), .B(n8735), .Z(n1899) );
  OR2 U4640 ( .A(n8728), .B(n8736), .Z(n1897) );
  OR2 U4641 ( .A(n5249), .B(n8737), .Z(n1896) );
  OR2 U4642 ( .A(n8738), .B(n8739), .Z(n1895) );
  OR2 U4643 ( .A(n5247), .B(n8728), .Z(n8739) );
  OR2 U4644 ( .A(n8740), .B(n8741), .Z(n1894) );
  OR2 U4645 ( .A(n8734), .B(n8742), .Z(n8741) );
  OR2 U4646 ( .A(n5254), .B(n8743), .Z(n8740) );
  OR2 U4647 ( .A(n8744), .B(n8745), .Z(n8743) );
  OR2 U4648 ( .A(n8738), .B(n8732), .Z(n1893) );
  OR2 U4649 ( .A(n5249), .B(n5248), .Z(n8732) );
  OR2 U4650 ( .A(n8746), .B(n8747), .Z(n1892) );
  OR2 U4651 ( .A(n8742), .B(n8748), .Z(n8747) );
  OR2 U4652 ( .A(n5257), .B(n8734), .Z(n8746) );
  OR2 U4653 ( .A(n8738), .B(n8749), .Z(n1891) );
  OR2 U4654 ( .A(n5248), .B(n8728), .Z(n8749) );
  OR2 U4655 ( .A(n8750), .B(n8751), .Z(n1890) );
  OR2 U4656 ( .A(n5254), .B(n8731), .Z(n8751) );
  OR2 U4657 ( .A(n8744), .B(n8752), .Z(n8750) );
  OR2 U4658 ( .A(n5257), .B(n8753), .Z(n8752) );
  OR2 U4659 ( .A(n8738), .B(n8754), .Z(n1889) );
  OR2 U4660 ( .A(n5249), .B(n5247), .Z(n8754) );
  OR2 U4661 ( .A(n8755), .B(n5245), .Z(n8738) );
  OR2 U4662 ( .A(n8756), .B(n8757), .Z(n1888) );
  OR2 U4663 ( .A(n8753), .B(n8745), .Z(n8756) );
  OR2 U4664 ( .A(n8734), .B(n8736), .Z(n1887) );
  OR2 U4665 ( .A(n8758), .B(n8759), .Z(n1886) );
  OR2 U4666 ( .A(n8731), .B(n8760), .Z(n8759) );
  OR2 U4667 ( .A(n8761), .B(n8762), .Z(n1885) );
  OR2 U4668 ( .A(n8763), .B(n8764), .Z(n8762) );
  OR2 U4669 ( .A(n8761), .B(n8765), .Z(n1884) );
  OR2 U4670 ( .A(n8766), .B(n8767), .Z(n8765) );
  OR2 U4671 ( .A(n8768), .B(n8769), .Z(n8761) );
  AN2 U4672 ( .A(n8770), .B(n5442), .Z(n8769) );
  AN2 U4673 ( .A(n8721), .B(n8771), .Z(n8768) );
  OR2 U4674 ( .A(n5444), .B(n5443), .Z(n8771) );
  IV U4675 ( .A(n1298), .Z(n5444) );
  OR2 U4676 ( .A(n8772), .B(n8773), .Z(n1883) );
  OR2 U4677 ( .A(n8774), .B(n8775), .Z(n8773) );
  OR2 U4678 ( .A(n8772), .B(n8776), .Z(n1882) );
  OR2 U4679 ( .A(n8777), .B(n8778), .Z(n8776) );
  OR2 U4680 ( .A(n8779), .B(n8780), .Z(n8772) );
  AN2 U4681 ( .A(n8781), .B(n5424), .Z(n8780) );
  AN2 U4682 ( .A(n8723), .B(n8782), .Z(n8779) );
  OR2 U4683 ( .A(n5426), .B(n5425), .Z(n8782) );
  IV U4684 ( .A(n1318), .Z(n5426) );
  OR2 U4685 ( .A(n8783), .B(n8784), .Z(n1881) );
  OR2 U4686 ( .A(n8785), .B(n8786), .Z(n8784) );
  OR2 U4687 ( .A(n8783), .B(n8787), .Z(n1880) );
  OR2 U4688 ( .A(n8788), .B(n8789), .Z(n8787) );
  OR2 U4689 ( .A(n8790), .B(n8791), .Z(n8783) );
  AN2 U4690 ( .A(n8792), .B(n5406), .Z(n8791) );
  AN2 U4691 ( .A(n8725), .B(n8793), .Z(n8790) );
  OR2 U4692 ( .A(n5408), .B(n5407), .Z(n8793) );
  IV U4693 ( .A(n1337), .Z(n5408) );
  OR2 U4694 ( .A(n8794), .B(n8795), .Z(n1879) );
  OR2 U4695 ( .A(n8796), .B(n8797), .Z(n8795) );
  OR2 U4696 ( .A(n8794), .B(n8798), .Z(n1878) );
  OR2 U4697 ( .A(n8799), .B(n8800), .Z(n8798) );
  OR2 U4698 ( .A(n8801), .B(n8802), .Z(n8794) );
  AN2 U4699 ( .A(n8803), .B(n5387), .Z(n8802) );
  AN2 U4700 ( .A(n8727), .B(n8804), .Z(n8801) );
  OR2 U4701 ( .A(n5389), .B(n5388), .Z(n8804) );
  IV U4702 ( .A(n1358), .Z(n5389) );
  OR2 U4703 ( .A(n8805), .B(n8806), .Z(n1877) );
  OR2 U4704 ( .A(n8807), .B(n8808), .Z(n8806) );
  OR2 U4705 ( .A(n8805), .B(n8809), .Z(n1876) );
  OR2 U4706 ( .A(n8810), .B(n8811), .Z(n8809) );
  OR2 U4707 ( .A(n8812), .B(n8813), .Z(n8805) );
  AN2 U4708 ( .A(n8814), .B(n5367), .Z(n8813) );
  IV U4709 ( .A(n1519), .Z(n5367) );
  AN2 U4710 ( .A(n8815), .B(n8816), .Z(n8812) );
  OR2 U4711 ( .A(n5369), .B(n5368), .Z(n8816) );
  IV U4712 ( .A(n1278), .Z(n5369) );
  OR2 U4713 ( .A(n8817), .B(n8818), .Z(n1875) );
  OR2 U4714 ( .A(n8819), .B(n8820), .Z(n8818) );
  OR2 U4715 ( .A(n8817), .B(n8821), .Z(n1874) );
  OR2 U4716 ( .A(n8822), .B(n8823), .Z(n8821) );
  OR2 U4717 ( .A(n8824), .B(n8825), .Z(n8817) );
  AN2 U4718 ( .A(n8826), .B(n5349), .Z(n8825) );
  AN2 U4719 ( .A(n8827), .B(n8828), .Z(n8824) );
  OR2 U4720 ( .A(n5351), .B(n5350), .Z(n8828) );
  IV U4721 ( .A(n1288), .Z(n5351) );
  OR2 U4722 ( .A(n8829), .B(n8830), .Z(n1873) );
  OR2 U4723 ( .A(n8831), .B(n8832), .Z(n8830) );
  OR2 U4724 ( .A(n8829), .B(n8833), .Z(n1872) );
  OR2 U4725 ( .A(n8834), .B(n8835), .Z(n8833) );
  OR2 U4726 ( .A(n8836), .B(n8837), .Z(n8829) );
  AN2 U4727 ( .A(n8838), .B(n5331), .Z(n8837) );
  AN2 U4728 ( .A(n8839), .B(n8840), .Z(n8836) );
  OR2 U4729 ( .A(n5333), .B(n5332), .Z(n8840) );
  IV U4730 ( .A(n1308), .Z(n5333) );
  OR2 U4731 ( .A(n8841), .B(n8842), .Z(n1871) );
  OR2 U4732 ( .A(n8843), .B(n8844), .Z(n8842) );
  OR2 U4733 ( .A(n8841), .B(n8845), .Z(n1870) );
  OR2 U4734 ( .A(n8846), .B(n8847), .Z(n8845) );
  OR2 U4735 ( .A(n8848), .B(n8849), .Z(n8841) );
  AN2 U4736 ( .A(n8850), .B(n5312), .Z(n8849) );
  AN2 U4737 ( .A(n8851), .B(n8852), .Z(n8848) );
  OR2 U4738 ( .A(n5314), .B(n5313), .Z(n8852) );
  IV U4739 ( .A(n1327), .Z(n5314) );
  AN2 U4740 ( .A(n8853), .B(n8815), .Z(n175) );
  AN2 U4741 ( .A(n1371), .B(n1278), .Z(n8853) );
  AN2 U4742 ( .A(n8854), .B(n8827), .Z(n159) );
  AN2 U4743 ( .A(n1384), .B(n1288), .Z(n8854) );
  AN2 U4744 ( .A(n8855), .B(n8839), .Z(n143) );
  AN2 U4745 ( .A(n1410), .B(n1308), .Z(n8855) );
  AN2 U4746 ( .A(n8856), .B(n8851), .Z(n127) );
  AN2 U4747 ( .A(n1433), .B(n1327), .Z(n8856) );
  AN2 U4748 ( .A(tx_fifo_pop_2), .B(n5684), .Z(n1115) );
  OR2 U4749 ( .A(n8857), .B(n8858), .Z(U8_Z_9) );
  OR2 U4750 ( .A(n8859), .B(n8860), .Z(n8858) );
  AN2 U4751 ( .A(n8861), .B(n8862), .Z(n8860) );
  IV U4752 ( .A(U3_U1_DATA3_9), .Z(n8862) );
  AN2 U4753 ( .A(U3_U1_DATA3_9), .B(n8863), .Z(n8859) );
  AN2 U4754 ( .A(n8864), .B(n8865), .Z(U8_Z_8) );
  OR2 U4755 ( .A(n8866), .B(n8861), .Z(n8865) );
  IV U4756 ( .A(n8863), .Z(n8861) );
  AN2 U4757 ( .A(U3_U1_DATA3_8), .B(n8867), .Z(n8866) );
  AN2 U4758 ( .A(n8864), .B(n8868), .Z(U8_Z_7) );
  OR2 U4759 ( .A(n8869), .B(n8870), .Z(n8868) );
  IV U4760 ( .A(n8867), .Z(n8870) );
  AN2 U4761 ( .A(U3_U1_DATA3_7), .B(n8871), .Z(n8869) );
  OR2 U4762 ( .A(n8857), .B(n8872), .Z(U8_Z_6) );
  OR2 U4763 ( .A(n8873), .B(n8874), .Z(n8872) );
  AN2 U4764 ( .A(U3_U1_DATA3_6), .B(n8875), .Z(n8874) );
  IV U4765 ( .A(n8871), .Z(n8873) );
  AN2 U4766 ( .A(n8864), .B(n8876), .Z(U8_Z_5) );
  OR2 U4767 ( .A(n8877), .B(n8878), .Z(n8876) );
  IV U4768 ( .A(n8875), .Z(n8878) );
  AN2 U4769 ( .A(U3_U1_DATA3_5), .B(n8879), .Z(n8877) );
  AN2 U4770 ( .A(n8864), .B(n8880), .Z(U8_Z_4) );
  OR2 U4771 ( .A(n8881), .B(n8882), .Z(n8880) );
  IV U4772 ( .A(n8879), .Z(n8882) );
  AN2 U4773 ( .A(U3_U1_DATA3_4), .B(n8883), .Z(n8881) );
  OR2 U4774 ( .A(n8857), .B(n8884), .Z(U8_Z_3) );
  OR2 U4775 ( .A(n8885), .B(n8886), .Z(n8884) );
  AN2 U4776 ( .A(U3_U1_DATA3_3), .B(n8887), .Z(n8886) );
  IV U4777 ( .A(n8883), .Z(n8885) );
  AN2 U4778 ( .A(n8864), .B(n8888), .Z(U8_Z_2) );
  OR2 U4779 ( .A(n8889), .B(n8890), .Z(n8888) );
  IV U4780 ( .A(n8887), .Z(n8890) );
  AN2 U4781 ( .A(U3_U1_DATA3_2), .B(n8891), .Z(n8889) );
  IV U4782 ( .A(n8857), .Z(n8864) );
  OR2 U4783 ( .A(n8857), .B(n8892), .Z(U8_Z_10) );
  OR2 U4784 ( .A(n8893), .B(n8894), .Z(n8892) );
  IV U4785 ( .A(n8895), .Z(n8894) );
  OR2 U4786 ( .A(n8896), .B(U3_U1_DATA3_10), .Z(n8895) );
  AN2 U4787 ( .A(U3_U1_DATA3_10), .B(n8896), .Z(n8893) );
  OR2 U4788 ( .A(U3_U1_DATA3_9), .B(n8863), .Z(n8896) );
  OR2 U4789 ( .A(U3_U1_DATA3_8), .B(n8867), .Z(n8863) );
  OR2 U4790 ( .A(U3_U1_DATA3_7), .B(n8871), .Z(n8867) );
  OR2 U4791 ( .A(U3_U1_DATA3_6), .B(n8875), .Z(n8871) );
  OR2 U4792 ( .A(U3_U1_DATA3_5), .B(n8879), .Z(n8875) );
  OR2 U4793 ( .A(U3_U1_DATA3_4), .B(n8883), .Z(n8879) );
  OR2 U4794 ( .A(U3_U1_DATA3_3), .B(n8887), .Z(n8883) );
  OR2 U4795 ( .A(U3_U1_DATA3_2), .B(n8891), .Z(n8887) );
  OR2 U4796 ( .A(n8857), .B(n8897), .Z(U8_Z_1) );
  OR2 U4797 ( .A(n8898), .B(n8899), .Z(n8897) );
  AN2 U4798 ( .A(U3_U1_DATA3_1), .B(n8900), .Z(n8899) );
  IV U4799 ( .A(n8891), .Z(n8898) );
  OR2 U4800 ( .A(U3_U1_DATA3_1), .B(n8900), .Z(n8891) );
  OR2 U4801 ( .A(n8857), .B(n8901), .Z(U8_Z_0) );
  OR2 U4802 ( .A(n8902), .B(n8903), .Z(n8901) );
  AN2 U4803 ( .A(U3_U1_DATA3_0), .B(n5538), .Z(n8903) );
  IV U4804 ( .A(n8900), .Z(n8902) );
  OR2 U4805 ( .A(U3_U1_DATA3_0), .B(n5538), .Z(n8900) );
  IV U4806 ( .A(sub_125_aco_B_0_), .Z(n5538) );
  OR2 U4807 ( .A(n8904), .B(n8905), .Z(U7_Z_9) );
  OR2 U4808 ( .A(n8906), .B(n8907), .Z(n8905) );
  AN2 U4809 ( .A(sub_126_aco_A_9_), .B(n8908), .Z(n8907) );
  IV U4810 ( .A(n8909), .Z(n8906) );
  AN2 U4811 ( .A(n8910), .B(n8911), .Z(U7_Z_8) );
  OR2 U4812 ( .A(n8912), .B(n8913), .Z(n8911) );
  IV U4813 ( .A(n8908), .Z(n8913) );
  AN2 U4814 ( .A(sub_126_aco_A_8_), .B(n8914), .Z(n8912) );
  OR2 U4815 ( .A(n8904), .B(n8915), .Z(U7_Z_7) );
  OR2 U4816 ( .A(n8916), .B(n8917), .Z(n8915) );
  AN2 U4817 ( .A(sub_126_aco_A_7_), .B(n8918), .Z(n8917) );
  IV U4818 ( .A(n8914), .Z(n8916) );
  OR2 U4819 ( .A(n8904), .B(n8919), .Z(U7_Z_6) );
  OR2 U4820 ( .A(n8920), .B(n8921), .Z(n8919) );
  AN2 U4821 ( .A(sub_126_aco_A_6_), .B(n8922), .Z(n8921) );
  IV U4822 ( .A(n8918), .Z(n8920) );
  OR2 U4823 ( .A(n8904), .B(n8923), .Z(U7_Z_5) );
  OR2 U4824 ( .A(n8924), .B(n8925), .Z(n8923) );
  AN2 U4825 ( .A(sub_126_aco_A_5_), .B(n8926), .Z(n8925) );
  IV U4826 ( .A(n8922), .Z(n8924) );
  OR2 U4827 ( .A(n8904), .B(n8927), .Z(U7_Z_4) );
  OR2 U4828 ( .A(n8928), .B(n8929), .Z(n8927) );
  AN2 U4829 ( .A(sub_126_aco_A_4_), .B(n8930), .Z(n8929) );
  IV U4830 ( .A(n8926), .Z(n8928) );
  OR2 U4831 ( .A(n8904), .B(n8931), .Z(U7_Z_3) );
  OR2 U4832 ( .A(n8932), .B(n8933), .Z(n8931) );
  AN2 U4833 ( .A(sub_126_aco_A_3_), .B(n8934), .Z(n8933) );
  IV U4834 ( .A(n8930), .Z(n8932) );
  AN2 U4835 ( .A(n8910), .B(n8935), .Z(U7_Z_2) );
  OR2 U4836 ( .A(n8936), .B(n8937), .Z(n8935) );
  IV U4837 ( .A(n8934), .Z(n8937) );
  AN2 U4838 ( .A(sub_126_aco_A_2_), .B(n8938), .Z(n8936) );
  OR2 U4839 ( .A(n8904), .B(n8939), .Z(U7_Z_19) );
  OR2 U4840 ( .A(n8940), .B(n8941), .Z(n8939) );
  IV U4841 ( .A(n8942), .Z(n8941) );
  OR2 U4842 ( .A(n8943), .B(sub_126_aco_A_19_), .Z(n8942) );
  AN2 U4843 ( .A(sub_126_aco_A_19_), .B(n8943), .Z(n8940) );
  OR2 U4844 ( .A(sub_126_aco_A_18_), .B(n8944), .Z(n8943) );
  AN2 U4845 ( .A(n8910), .B(n8945), .Z(U7_Z_18) );
  OR2 U4846 ( .A(n8946), .B(n8947), .Z(n8945) );
  AN2 U4847 ( .A(n8948), .B(n8949), .Z(n8947) );
  IV U4848 ( .A(sub_126_aco_A_18_), .Z(n8949) );
  AN2 U4849 ( .A(sub_126_aco_A_18_), .B(n8944), .Z(n8946) );
  AN2 U4850 ( .A(n8910), .B(n8950), .Z(U7_Z_17) );
  OR2 U4851 ( .A(n8951), .B(n8948), .Z(n8950) );
  IV U4852 ( .A(n8944), .Z(n8948) );
  OR2 U4853 ( .A(sub_126_aco_A_17_), .B(n8952), .Z(n8944) );
  AN2 U4854 ( .A(sub_126_aco_A_17_), .B(n8952), .Z(n8951) );
  AN2 U4855 ( .A(n8910), .B(n8953), .Z(U7_Z_16) );
  OR2 U4856 ( .A(n8954), .B(n8955), .Z(n8953) );
  IV U4857 ( .A(n8952), .Z(n8955) );
  OR2 U4858 ( .A(sub_126_aco_A_16_), .B(n8956), .Z(n8952) );
  AN2 U4859 ( .A(sub_126_aco_A_16_), .B(n8956), .Z(n8954) );
  OR2 U4860 ( .A(n8904), .B(n8957), .Z(U7_Z_15) );
  OR2 U4861 ( .A(n8958), .B(n8959), .Z(n8957) );
  AN2 U4862 ( .A(sub_126_aco_A_15_), .B(n8960), .Z(n8959) );
  IV U4863 ( .A(n8956), .Z(n8958) );
  OR2 U4864 ( .A(sub_126_aco_A_15_), .B(n8960), .Z(n8956) );
  AN2 U4865 ( .A(n8910), .B(n8961), .Z(U7_Z_14) );
  OR2 U4866 ( .A(n8962), .B(n8963), .Z(n8961) );
  IV U4867 ( .A(n8960), .Z(n8963) );
  OR2 U4868 ( .A(sub_126_aco_A_14_), .B(n8964), .Z(n8960) );
  AN2 U4869 ( .A(sub_126_aco_A_14_), .B(n8964), .Z(n8962) );
  AN2 U4870 ( .A(n8910), .B(n8965), .Z(U7_Z_13) );
  OR2 U4871 ( .A(n8966), .B(n8967), .Z(n8965) );
  IV U4872 ( .A(n8964), .Z(n8967) );
  OR2 U4873 ( .A(sub_126_aco_A_13_), .B(n8968), .Z(n8964) );
  AN2 U4874 ( .A(sub_126_aco_A_13_), .B(n8968), .Z(n8966) );
  OR2 U4875 ( .A(n8904), .B(n8969), .Z(U7_Z_12) );
  OR2 U4876 ( .A(n8970), .B(n8971), .Z(n8969) );
  AN2 U4877 ( .A(sub_126_aco_A_12_), .B(n8972), .Z(n8971) );
  IV U4878 ( .A(n8968), .Z(n8970) );
  OR2 U4879 ( .A(sub_126_aco_A_12_), .B(n8972), .Z(n8968) );
  OR2 U4880 ( .A(n8904), .B(n8973), .Z(U7_Z_11) );
  OR2 U4881 ( .A(n8974), .B(n8975), .Z(n8973) );
  AN2 U4882 ( .A(sub_126_aco_A_11_), .B(n8976), .Z(n8975) );
  IV U4883 ( .A(n8972), .Z(n8974) );
  OR2 U4884 ( .A(sub_126_aco_A_11_), .B(n8976), .Z(n8972) );
  AN2 U4885 ( .A(n8910), .B(n8977), .Z(U7_Z_10) );
  OR2 U4886 ( .A(n8978), .B(n8979), .Z(n8977) );
  IV U4887 ( .A(n8976), .Z(n8979) );
  OR2 U4888 ( .A(sub_126_aco_A_10_), .B(n8909), .Z(n8976) );
  AN2 U4889 ( .A(sub_126_aco_A_10_), .B(n8909), .Z(n8978) );
  OR2 U4890 ( .A(sub_126_aco_A_9_), .B(n8908), .Z(n8909) );
  OR2 U4891 ( .A(sub_126_aco_A_8_), .B(n8914), .Z(n8908) );
  OR2 U4892 ( .A(sub_126_aco_A_7_), .B(n8918), .Z(n8914) );
  OR2 U4893 ( .A(sub_126_aco_A_6_), .B(n8922), .Z(n8918) );
  OR2 U4894 ( .A(sub_126_aco_A_5_), .B(n8926), .Z(n8922) );
  OR2 U4895 ( .A(sub_126_aco_A_4_), .B(n8930), .Z(n8926) );
  OR2 U4896 ( .A(sub_126_aco_A_3_), .B(n8934), .Z(n8930) );
  OR2 U4897 ( .A(sub_126_aco_A_2_), .B(n8938), .Z(n8934) );
  IV U4898 ( .A(n8904), .Z(n8910) );
  OR2 U4899 ( .A(n8904), .B(n8980), .Z(U7_Z_1) );
  OR2 U4900 ( .A(n8981), .B(n8982), .Z(n8980) );
  AN2 U4901 ( .A(sub_126_aco_A_1_), .B(n8983), .Z(n8982) );
  IV U4902 ( .A(n8938), .Z(n8981) );
  OR2 U4903 ( .A(sub_126_aco_A_1_), .B(n8983), .Z(n8938) );
  OR2 U4904 ( .A(n8904), .B(n8984), .Z(U7_Z_0) );
  OR2 U4905 ( .A(n8985), .B(n8986), .Z(n8984) );
  AN2 U4906 ( .A(sub_126_aco_A_0_), .B(n5559), .Z(n8986) );
  IV U4907 ( .A(n8983), .Z(n8985) );
  OR2 U4908 ( .A(sub_126_aco_A_0_), .B(n5559), .Z(n8983) );
  IV U4909 ( .A(sub_126_aco_B_0_), .Z(n5559) );
  AN2 U4910 ( .A(n2664), .B(n8987), .Z(U67_Z_3) );
  OR2 U4911 ( .A(n8988), .B(n8989), .Z(n8987) );
  OR2 U4912 ( .A(n8904), .B(n8990), .Z(n8989) );
  OR2 U4913 ( .A(n8991), .B(n8857), .Z(n8988) );
  OR2 U4914 ( .A(n8992), .B(n8993), .Z(n8857) );
  AN2 U4915 ( .A(U76_DATA3_0), .B(n8717), .Z(n8992) );
  AN2 U4916 ( .A(n8994), .B(U111_DATA3_0), .Z(n8991) );
  AN2 U4917 ( .A(n2664), .B(n8995), .Z(U67_Z_2) );
  OR2 U4918 ( .A(n8996), .B(n8997), .Z(n8995) );
  OR2 U4919 ( .A(n8998), .B(n8990), .Z(n8997) );
  OR2 U4920 ( .A(n8999), .B(n9000), .Z(n8990) );
  AN2 U4921 ( .A(n8994), .B(U112_DATA3_0), .Z(n8998) );
  OR2 U4922 ( .A(n9001), .B(n9002), .Z(n8994) );
  OR2 U4923 ( .A(n9003), .B(n8715), .Z(n9002) );
  OR2 U4924 ( .A(n9004), .B(n9005), .Z(n8996) );
  AN2 U4925 ( .A(n2664), .B(n9006), .Z(U67_Z_1) );
  OR2 U4926 ( .A(n9007), .B(n9008), .Z(n9006) );
  OR2 U4927 ( .A(n9009), .B(n9010), .Z(n9008) );
  AN2 U4928 ( .A(n2753), .B(n8662), .Z(n9009) );
  OR2 U4929 ( .A(n9011), .B(n9012), .Z(n9007) );
  AN2 U4930 ( .A(n9013), .B(U113_DATA3_0), .Z(n9012) );
  AN2 U4931 ( .A(n2664), .B(n9014), .Z(U67_Z_0) );
  OR2 U4932 ( .A(n9015), .B(n9016), .Z(n9014) );
  OR2 U4933 ( .A(n8993), .B(n9010), .Z(n9016) );
  OR2 U4934 ( .A(n9017), .B(n9018), .Z(n9010) );
  AN2 U4935 ( .A(n2770), .B(n8719), .Z(n9018) );
  OR2 U4936 ( .A(n9019), .B(n9020), .Z(n8993) );
  AN2 U4937 ( .A(U76_DATA4_0), .B(n5482), .Z(n9019) );
  OR2 U4938 ( .A(n9021), .B(n9022), .Z(n9015) );
  AN2 U4939 ( .A(n2762), .B(n8717), .Z(n9022) );
  AN2 U4940 ( .A(n9013), .B(U114_DATA2_0), .Z(n9021) );
  OR2 U4941 ( .A(n9001), .B(n9023), .Z(n9013) );
  OR2 U4942 ( .A(n9024), .B(n9025), .Z(n9023) );
  OR2 U4943 ( .A(n9026), .B(n9027), .Z(n9001) );
  OR2 U4944 ( .A(n9028), .B(n9029), .Z(n9027) );
  AN2 U4945 ( .A(n4903), .B(n8719), .Z(n9029) );
  IV U4946 ( .A(n9030), .Z(n4903) );
  OR2 U4947 ( .A(U71_DATA3_0), .B(U69_DATA2_0), .Z(n9030) );
  AN2 U4948 ( .A(n2664), .B(n9031), .Z(U66_Z_1) );
  OR2 U4949 ( .A(n9032), .B(n9033), .Z(n9031) );
  AN2 U4950 ( .A(n9034), .B(tx_mode[1]), .Z(n9032) );
  OR2 U4951 ( .A(n9035), .B(n8661), .Z(n9034) );
  AN2 U4952 ( .A(n2664), .B(n9036), .Z(U66_Z_0) );
  OR2 U4953 ( .A(n9037), .B(n8904), .Z(n9036) );
  OR2 U4954 ( .A(n9038), .B(n9011), .Z(n8904) );
  AN2 U4955 ( .A(n9039), .B(tx_mode[0]), .Z(n9037) );
  OR2 U4956 ( .A(n9035), .B(n9040), .Z(n9039) );
  OR2 U4957 ( .A(n9003), .B(n9041), .Z(n9040) );
  IV U4958 ( .A(n9042), .Z(n9041) );
  OR2 U4959 ( .A(n9043), .B(U69_DATA2_0), .Z(n9042) );
  OR2 U4960 ( .A(n9044), .B(n9045), .Z(n9035) );
  OR2 U4961 ( .A(n9046), .B(n9047), .Z(n9045) );
  AN2 U4962 ( .A(n2756), .B(n8662), .Z(n9046) );
  OR2 U4963 ( .A(n9025), .B(n9048), .Z(n9044) );
  OR2 U4964 ( .A(n9028), .B(n9049), .Z(n9048) );
  AN2 U4965 ( .A(n2747), .B(n5482), .Z(n9049) );
  AN2 U4966 ( .A(n9050), .B(n4898), .Z(n9028) );
  IV U4967 ( .A(n9051), .Z(n4898) );
  OR2 U4968 ( .A(n3273), .B(U72_DATA3_0), .Z(n9051) );
  AN2 U4969 ( .A(n8715), .B(sub_128_aco_B_0_), .Z(n9025) );
  AN2 U4970 ( .A(n2664), .B(n9052), .Z(U65_Z_0) );
  OR2 U4971 ( .A(n9053), .B(n9004), .Z(n9052) );
  AN2 U4972 ( .A(U107_DATA1_0), .B(n9054), .Z(n9053) );
  OR2 U4973 ( .A(n9055), .B(n9056), .Z(n9054) );
  OR2 U4974 ( .A(n8661), .B(n9057), .Z(n9056) );
  OR2 U4975 ( .A(n9026), .B(n9058), .Z(n9055) );
  OR2 U4976 ( .A(n9005), .B(n9038), .Z(n9058) );
  AN2 U4977 ( .A(U72_DATA2_0), .B(n8662), .Z(n9038) );
  OR2 U4978 ( .A(n9059), .B(n9060), .Z(n9026) );
  OR2 U4979 ( .A(n9061), .B(n9062), .Z(n9060) );
  AN2 U4980 ( .A(n4894), .B(n5482), .Z(n9062) );
  IV U4981 ( .A(n9063), .Z(n4894) );
  OR2 U4982 ( .A(U76_DATA4_0), .B(U73_DATA6_0), .Z(n9063) );
  AN2 U4983 ( .A(n9064), .B(n9065), .Z(n9061) );
  AN2 U4984 ( .A(n9066), .B(n9067), .Z(n9065) );
  IV U4985 ( .A(U76_DATA3_0), .Z(n9067) );
  IV U4986 ( .A(n9068), .Z(n9064) );
  OR2 U4987 ( .A(n9069), .B(U69_DATA4_0), .Z(n9068) );
  AN2 U4988 ( .A(n4899), .B(n8662), .Z(n9059) );
  IV U4989 ( .A(n9070), .Z(n4899) );
  OR2 U4990 ( .A(U72_DATA2_0), .B(n9071), .Z(n9070) );
  OR2 U4991 ( .A(n3273), .B(n2593), .Z(n9071) );
  AN2 U4992 ( .A(n2664), .B(n9072), .Z(U64_Z_0) );
  OR2 U4993 ( .A(n9073), .B(n9005), .Z(n9072) );
  AN2 U4994 ( .A(n8662), .B(n2593), .Z(n9005) );
  AN2 U4995 ( .A(TXxREFRESH), .B(n9074), .Z(n9073) );
  OR2 U4996 ( .A(n9075), .B(n9076), .Z(n9074) );
  OR2 U4997 ( .A(n9057), .B(n9077), .Z(n9076) );
  OR2 U4998 ( .A(n9078), .B(n9047), .Z(n9077) );
  OR2 U4999 ( .A(n9079), .B(n9080), .Z(n9047) );
  OR2 U5000 ( .A(n9004), .B(n9020), .Z(n9080) );
  AN2 U5001 ( .A(n2534), .B(n9081), .Z(n9020) );
  AN2 U5002 ( .A(n4900), .B(n2533), .Z(n9081) );
  AN2 U5003 ( .A(n8717), .B(n9082), .Z(n9079) );
  OR2 U5004 ( .A(U76_DATA3_0), .B(n9066), .Z(n9082) );
  IV U5005 ( .A(U73_DATA5_0), .Z(n9066) );
  AN2 U5006 ( .A(n2771), .B(n8719), .Z(n9078) );
  OR2 U5007 ( .A(n9083), .B(n8715), .Z(n9057) );
  IV U5008 ( .A(n9084), .Z(n8715) );
  AN2 U5009 ( .A(n9050), .B(n4900), .Z(n9083) );
  IV U5010 ( .A(n3273), .Z(n4900) );
  OR2 U5011 ( .A(n9085), .B(n9086), .Z(n9075) );
  OR2 U5012 ( .A(n5482), .B(n9087), .Z(n9086) );
  AN2 U5013 ( .A(n2757), .B(n8662), .Z(n9087) );
  IV U5014 ( .A(n9088), .Z(n5482) );
  OR2 U5015 ( .A(n2559), .B(n2560), .Z(n9088) );
  OR2 U5016 ( .A(n2587), .B(n9024), .Z(n9085) );
  AN2 U5017 ( .A(n2664), .B(n9089), .Z(U63_Z_0) );
  OR2 U5018 ( .A(n9090), .B(n9011), .Z(n9089) );
  AN2 U5019 ( .A(TXxQUIET), .B(n9091), .Z(n9090) );
  OR2 U5020 ( .A(n9092), .B(n9093), .Z(n9091) );
  OR2 U5021 ( .A(n2775), .B(n9003), .Z(n9093) );
  AN2 U5022 ( .A(n9094), .B(n9024), .Z(n9003) );
  IV U5023 ( .A(n2517), .Z(n9094) );
  AN2 U5024 ( .A(n2749), .B(n9050), .Z(n9092) );
  AN2 U5025 ( .A(n9095), .B(n9096), .Z(U6_Z_9) );
  OR2 U5026 ( .A(n9097), .B(n9098), .Z(n9095) );
  AN2 U5027 ( .A(sub_127_aco_A_9_), .B(n9099), .Z(n9097) );
  OR2 U5028 ( .A(n9100), .B(n9101), .Z(U6_Z_8) );
  OR2 U5029 ( .A(n9000), .B(n9102), .Z(n9101) );
  IV U5030 ( .A(n9099), .Z(n9102) );
  AN2 U5031 ( .A(sub_127_aco_A_8_), .B(n9103), .Z(n9100) );
  OR2 U5032 ( .A(n9104), .B(n9105), .Z(U6_Z_7) );
  OR2 U5033 ( .A(n9000), .B(n9106), .Z(n9105) );
  IV U5034 ( .A(n9103), .Z(n9106) );
  AN2 U5035 ( .A(sub_127_aco_A_7_), .B(n9107), .Z(n9104) );
  OR2 U5036 ( .A(n9108), .B(n9109), .Z(U6_Z_6) );
  OR2 U5037 ( .A(n9000), .B(n9110), .Z(n9109) );
  IV U5038 ( .A(n9107), .Z(n9110) );
  AN2 U5039 ( .A(sub_127_aco_A_6_), .B(n9111), .Z(n9108) );
  AN2 U5040 ( .A(n9112), .B(n9096), .Z(U6_Z_5) );
  OR2 U5041 ( .A(n9113), .B(n9114), .Z(n9112) );
  IV U5042 ( .A(n9111), .Z(n9114) );
  AN2 U5043 ( .A(sub_127_aco_A_5_), .B(n9115), .Z(n9113) );
  OR2 U5044 ( .A(n9116), .B(n9117), .Z(U6_Z_4) );
  OR2 U5045 ( .A(n9000), .B(n9118), .Z(n9117) );
  IV U5046 ( .A(n9115), .Z(n9118) );
  AN2 U5047 ( .A(sub_127_aco_A_4_), .B(n9119), .Z(n9116) );
  AN2 U5048 ( .A(n9120), .B(n9096), .Z(U6_Z_3) );
  OR2 U5049 ( .A(n9121), .B(n9122), .Z(n9120) );
  IV U5050 ( .A(n9119), .Z(n9122) );
  AN2 U5051 ( .A(sub_127_aco_A_3_), .B(n9123), .Z(n9121) );
  OR2 U5052 ( .A(n9124), .B(n9125), .Z(U6_Z_2) );
  OR2 U5053 ( .A(n9000), .B(n9126), .Z(n9125) );
  IV U5054 ( .A(n9123), .Z(n9126) );
  AN2 U5055 ( .A(sub_127_aco_A_2_), .B(n9127), .Z(n9124) );
  OR2 U5056 ( .A(n9000), .B(n9128), .Z(U6_Z_11) );
  OR2 U5057 ( .A(n9129), .B(n9130), .Z(n9128) );
  IV U5058 ( .A(n9131), .Z(n9130) );
  OR2 U5059 ( .A(n9132), .B(sub_127_aco_A_11_), .Z(n9131) );
  AN2 U5060 ( .A(sub_127_aco_A_11_), .B(n9132), .Z(n9129) );
  OR2 U5061 ( .A(sub_127_aco_A_10_), .B(n9133), .Z(n9132) );
  OR2 U5062 ( .A(n9000), .B(n9134), .Z(U6_Z_10) );
  OR2 U5063 ( .A(n9135), .B(n9136), .Z(n9134) );
  AN2 U5064 ( .A(n9098), .B(n9137), .Z(n9136) );
  IV U5065 ( .A(sub_127_aco_A_10_), .Z(n9137) );
  IV U5066 ( .A(n9133), .Z(n9098) );
  AN2 U5067 ( .A(sub_127_aco_A_10_), .B(n9133), .Z(n9135) );
  OR2 U5068 ( .A(sub_127_aco_A_9_), .B(n9099), .Z(n9133) );
  OR2 U5069 ( .A(sub_127_aco_A_8_), .B(n9103), .Z(n9099) );
  OR2 U5070 ( .A(sub_127_aco_A_7_), .B(n9107), .Z(n9103) );
  OR2 U5071 ( .A(sub_127_aco_A_6_), .B(n9111), .Z(n9107) );
  OR2 U5072 ( .A(sub_127_aco_A_5_), .B(n9115), .Z(n9111) );
  OR2 U5073 ( .A(sub_127_aco_A_4_), .B(n9119), .Z(n9115) );
  OR2 U5074 ( .A(sub_127_aco_A_3_), .B(n9123), .Z(n9119) );
  OR2 U5075 ( .A(sub_127_aco_A_2_), .B(n9127), .Z(n9123) );
  OR2 U5076 ( .A(n9138), .B(n9139), .Z(U6_Z_1) );
  OR2 U5077 ( .A(n9000), .B(n9140), .Z(n9139) );
  IV U5078 ( .A(n9127), .Z(n9140) );
  OR2 U5079 ( .A(sub_127_aco_A_1_), .B(n9141), .Z(n9127) );
  AN2 U5080 ( .A(sub_127_aco_A_1_), .B(n9141), .Z(n9138) );
  OR2 U5081 ( .A(n9142), .B(n9143), .Z(U6_Z_0) );
  OR2 U5082 ( .A(n9000), .B(n9144), .Z(n9143) );
  IV U5083 ( .A(n9141), .Z(n9144) );
  OR2 U5084 ( .A(sub_127_aco_A_0_), .B(n5572), .Z(n9141) );
  IV U5085 ( .A(n9096), .Z(n9000) );
  OR2 U5086 ( .A(sub_128_aco_B_0_), .B(n9084), .Z(n9096) );
  OR2 U5087 ( .A(n2551), .B(n2552), .Z(n9084) );
  AN2 U5088 ( .A(sub_127_aco_A_0_), .B(n5572), .Z(n9142) );
  IV U5089 ( .A(sub_127_aco_B_0_), .Z(n5572) );
  OR2 U5090 ( .A(n9145), .B(n9146), .Z(U5_Z_8) );
  OR2 U5091 ( .A(n9147), .B(n9148), .Z(n9146) );
  IV U5092 ( .A(n9149), .Z(n9148) );
  OR2 U5093 ( .A(n9150), .B(sub_128_aco_A_8_), .Z(n9149) );
  AN2 U5094 ( .A(sub_128_aco_A_8_), .B(n9150), .Z(n9147) );
  OR2 U5095 ( .A(sub_128_aco_A_7_), .B(n9151), .Z(n9150) );
  OR2 U5096 ( .A(n9145), .B(n9152), .Z(U5_Z_7) );
  OR2 U5097 ( .A(n9153), .B(n9154), .Z(n9152) );
  AN2 U5098 ( .A(n9155), .B(n9156), .Z(n9154) );
  IV U5099 ( .A(sub_128_aco_A_7_), .Z(n9156) );
  AN2 U5100 ( .A(sub_128_aco_A_7_), .B(n9151), .Z(n9153) );
  AN2 U5101 ( .A(n9157), .B(n9158), .Z(U5_Z_6) );
  OR2 U5102 ( .A(n9159), .B(n9155), .Z(n9158) );
  IV U5103 ( .A(n9151), .Z(n9155) );
  OR2 U5104 ( .A(sub_128_aco_A_6_), .B(n9160), .Z(n9151) );
  AN2 U5105 ( .A(sub_128_aco_A_6_), .B(n9160), .Z(n9159) );
  AN2 U5106 ( .A(n9157), .B(n9161), .Z(U5_Z_5) );
  OR2 U5107 ( .A(n9162), .B(n9163), .Z(n9161) );
  IV U5108 ( .A(n9160), .Z(n9163) );
  OR2 U5109 ( .A(sub_128_aco_A_5_), .B(n9164), .Z(n9160) );
  AN2 U5110 ( .A(sub_128_aco_A_5_), .B(n9164), .Z(n9162) );
  AN2 U5111 ( .A(n9157), .B(n9165), .Z(U5_Z_4) );
  OR2 U5112 ( .A(n9166), .B(n9167), .Z(n9165) );
  IV U5113 ( .A(n9164), .Z(n9167) );
  OR2 U5114 ( .A(sub_128_aco_A_4_), .B(n9168), .Z(n9164) );
  AN2 U5115 ( .A(sub_128_aco_A_4_), .B(n9168), .Z(n9166) );
  AN2 U5116 ( .A(n9157), .B(n9169), .Z(U5_Z_3) );
  OR2 U5117 ( .A(n9170), .B(n9171), .Z(n9169) );
  IV U5118 ( .A(n9168), .Z(n9171) );
  OR2 U5119 ( .A(sub_128_aco_A_3_), .B(n9172), .Z(n9168) );
  AN2 U5120 ( .A(sub_128_aco_A_3_), .B(n9172), .Z(n9170) );
  AN2 U5121 ( .A(n9157), .B(n9173), .Z(U5_Z_2) );
  OR2 U5122 ( .A(n9174), .B(n9175), .Z(n9173) );
  IV U5123 ( .A(n9172), .Z(n9175) );
  OR2 U5124 ( .A(sub_128_aco_A_2_), .B(n9176), .Z(n9172) );
  AN2 U5125 ( .A(sub_128_aco_A_2_), .B(n9176), .Z(n9174) );
  AN2 U5126 ( .A(n9157), .B(n9177), .Z(U5_Z_1) );
  OR2 U5127 ( .A(n9178), .B(n9179), .Z(n9177) );
  IV U5128 ( .A(n9176), .Z(n9179) );
  OR2 U5129 ( .A(sub_128_aco_A_1_), .B(n9180), .Z(n9176) );
  AN2 U5130 ( .A(sub_128_aco_A_1_), .B(n9180), .Z(n9178) );
  IV U5131 ( .A(n9145), .Z(n9157) );
  OR2 U5132 ( .A(n9145), .B(n9181), .Z(U5_Z_0) );
  OR2 U5133 ( .A(n9182), .B(n9183), .Z(n9181) );
  AN2 U5134 ( .A(sub_128_aco_A_0_), .B(n5582), .Z(n9183) );
  IV U5135 ( .A(n9180), .Z(n9182) );
  OR2 U5136 ( .A(sub_128_aco_A_0_), .B(n5582), .Z(n9180) );
  IV U5137 ( .A(sub_128_aco_B_0_), .Z(n5582) );
  OR2 U5138 ( .A(n9004), .B(n9033), .Z(n9145) );
  OR2 U5139 ( .A(n9017), .B(n9184), .Z(n9033) );
  AN2 U5140 ( .A(U69_DATA2_0), .B(n8719), .Z(n9184) );
  AN2 U5141 ( .A(n2517), .B(n9024), .Z(n9017) );
  AN2 U5142 ( .A(n8717), .B(U69_DATA4_0), .Z(n9004) );
  IV U5143 ( .A(n9069), .Z(n8717) );
  OR2 U5144 ( .A(n2555), .B(n2556), .Z(n9069) );
  OR2 U5145 ( .A(n9185), .B(n9186), .Z(U35_Z_9) );
  OR2 U5146 ( .A(n9187), .B(n9188), .Z(n9186) );
  OR2 U5147 ( .A(n9189), .B(n9190), .Z(n9188) );
  AN2 U5148 ( .A(U37_DATA4_9), .B(n9191), .Z(n9190) );
  AN2 U5149 ( .A(U37_DATA6_9), .B(n9192), .Z(n9189) );
  AN2 U5150 ( .A(U37_DATA1_9), .B(n9193), .Z(n9187) );
  OR2 U5151 ( .A(n9194), .B(n9195), .Z(n9185) );
  OR2 U5152 ( .A(n9196), .B(n9197), .Z(n9195) );
  AN2 U5153 ( .A(test_pat_seed_a[9]), .B(n9198), .Z(n9197) );
  AN2 U5154 ( .A(n9199), .B(n9200), .Z(n9196) );
  AN2 U5155 ( .A(test_pat_seed_b[9]), .B(n9201), .Z(n9194) );
  OR2 U5156 ( .A(n9202), .B(n9203), .Z(U35_Z_8) );
  OR2 U5157 ( .A(n9204), .B(n9205), .Z(n9203) );
  OR2 U5158 ( .A(n9206), .B(n9207), .Z(n9205) );
  AN2 U5159 ( .A(U37_DATA4_8), .B(n9191), .Z(n9207) );
  AN2 U5160 ( .A(U37_DATA6_8), .B(n9192), .Z(n9206) );
  AN2 U5161 ( .A(U37_DATA1_8), .B(n9193), .Z(n9204) );
  OR2 U5162 ( .A(n9208), .B(n9209), .Z(n9202) );
  OR2 U5163 ( .A(n9210), .B(n9211), .Z(n9209) );
  AN2 U5164 ( .A(test_pat_seed_a[8]), .B(n9198), .Z(n9211) );
  AN2 U5165 ( .A(n9199), .B(n9212), .Z(n9210) );
  AN2 U5166 ( .A(test_pat_seed_b[8]), .B(n9201), .Z(n9208) );
  OR2 U5167 ( .A(n9213), .B(n9214), .Z(U35_Z_7) );
  OR2 U5168 ( .A(n9215), .B(n9216), .Z(n9214) );
  OR2 U5169 ( .A(n9217), .B(n9218), .Z(n9216) );
  AN2 U5170 ( .A(U37_DATA4_7), .B(n9191), .Z(n9218) );
  AN2 U5171 ( .A(U37_DATA6_7), .B(n9192), .Z(n9217) );
  AN2 U5172 ( .A(U37_DATA1_7), .B(n9193), .Z(n9215) );
  OR2 U5173 ( .A(n9219), .B(n9220), .Z(n9213) );
  OR2 U5174 ( .A(n9221), .B(n9222), .Z(n9220) );
  AN2 U5175 ( .A(test_pat_seed_a[7]), .B(n9198), .Z(n9222) );
  AN2 U5176 ( .A(n9199), .B(n9223), .Z(n9221) );
  AN2 U5177 ( .A(test_pat_seed_b[7]), .B(n9201), .Z(n9219) );
  OR2 U5178 ( .A(n9224), .B(n9225), .Z(U35_Z_6) );
  OR2 U5179 ( .A(n9226), .B(n9227), .Z(n9225) );
  OR2 U5180 ( .A(n9228), .B(n9229), .Z(n9227) );
  AN2 U5181 ( .A(U37_DATA4_6), .B(n9191), .Z(n9229) );
  AN2 U5182 ( .A(U37_DATA6_6), .B(n9192), .Z(n9228) );
  AN2 U5183 ( .A(U37_DATA1_6), .B(n9193), .Z(n9226) );
  OR2 U5184 ( .A(n9230), .B(n9231), .Z(n9224) );
  OR2 U5185 ( .A(n9232), .B(n9233), .Z(n9231) );
  AN2 U5186 ( .A(test_pat_seed_a[6]), .B(n9198), .Z(n9233) );
  AN2 U5187 ( .A(n9234), .B(n9199), .Z(n9232) );
  AN2 U5188 ( .A(test_pat_seed_b[6]), .B(n9201), .Z(n9230) );
  OR2 U5189 ( .A(n9235), .B(n9236), .Z(U35_Z_57) );
  OR2 U5190 ( .A(n9237), .B(n9238), .Z(n9236) );
  OR2 U5191 ( .A(n9239), .B(n9240), .Z(n9238) );
  AN2 U5192 ( .A(U37_DATA4_57), .B(n9191), .Z(n9240) );
  AN2 U5193 ( .A(U37_DATA6_57), .B(n9192), .Z(n9239) );
  AN2 U5194 ( .A(U37_DATA1_57), .B(n9193), .Z(n9237) );
  OR2 U5195 ( .A(n9241), .B(n9242), .Z(n9235) );
  OR2 U5196 ( .A(n9243), .B(n9244), .Z(n9242) );
  AN2 U5197 ( .A(test_pat_seed_a[57]), .B(n9198), .Z(n9244) );
  AN2 U5198 ( .A(n9245), .B(n9199), .Z(n9243) );
  AN2 U5199 ( .A(test_pat_seed_b[57]), .B(n9201), .Z(n9241) );
  OR2 U5200 ( .A(n9246), .B(n9247), .Z(U35_Z_56) );
  OR2 U5201 ( .A(n9248), .B(n9249), .Z(n9247) );
  OR2 U5202 ( .A(n9250), .B(n9251), .Z(n9249) );
  AN2 U5203 ( .A(U37_DATA4_56), .B(n9191), .Z(n9251) );
  AN2 U5204 ( .A(U37_DATA6_56), .B(n9192), .Z(n9250) );
  AN2 U5205 ( .A(U37_DATA1_56), .B(n9193), .Z(n9248) );
  OR2 U5206 ( .A(n9252), .B(n9253), .Z(n9246) );
  OR2 U5207 ( .A(n9254), .B(n9255), .Z(n9253) );
  AN2 U5208 ( .A(test_pat_seed_a[56]), .B(n9198), .Z(n9255) );
  AN2 U5209 ( .A(n9256), .B(n9199), .Z(n9254) );
  AN2 U5210 ( .A(test_pat_seed_b[56]), .B(n9201), .Z(n9252) );
  OR2 U5211 ( .A(n9257), .B(n9258), .Z(U35_Z_55) );
  OR2 U5212 ( .A(n9259), .B(n9260), .Z(n9258) );
  OR2 U5213 ( .A(n9261), .B(n9262), .Z(n9260) );
  AN2 U5214 ( .A(U37_DATA4_55), .B(n9191), .Z(n9262) );
  AN2 U5215 ( .A(U37_DATA6_55), .B(n9192), .Z(n9261) );
  AN2 U5216 ( .A(U37_DATA1_55), .B(n9193), .Z(n9259) );
  OR2 U5217 ( .A(n9263), .B(n9264), .Z(n9257) );
  OR2 U5218 ( .A(n9265), .B(n9266), .Z(n9264) );
  AN2 U5219 ( .A(test_pat_seed_a[55]), .B(n9198), .Z(n9266) );
  AN2 U5220 ( .A(n9267), .B(n9199), .Z(n9265) );
  AN2 U5221 ( .A(test_pat_seed_b[55]), .B(n9201), .Z(n9263) );
  OR2 U5222 ( .A(n9268), .B(n9269), .Z(U35_Z_54) );
  OR2 U5223 ( .A(n9270), .B(n9271), .Z(n9269) );
  OR2 U5224 ( .A(n9272), .B(n9273), .Z(n9271) );
  AN2 U5225 ( .A(U37_DATA4_54), .B(n9191), .Z(n9273) );
  AN2 U5226 ( .A(U37_DATA6_54), .B(n9192), .Z(n9272) );
  AN2 U5227 ( .A(U37_DATA1_54), .B(n9193), .Z(n9270) );
  OR2 U5228 ( .A(n9274), .B(n9275), .Z(n9268) );
  OR2 U5229 ( .A(n9276), .B(n9277), .Z(n9275) );
  AN2 U5230 ( .A(test_pat_seed_a[54]), .B(n9198), .Z(n9277) );
  AN2 U5231 ( .A(n9278), .B(n9199), .Z(n9276) );
  AN2 U5232 ( .A(test_pat_seed_b[54]), .B(n9201), .Z(n9274) );
  OR2 U5233 ( .A(n9279), .B(n9280), .Z(U35_Z_53) );
  OR2 U5234 ( .A(n9281), .B(n9282), .Z(n9280) );
  OR2 U5235 ( .A(n9283), .B(n9284), .Z(n9282) );
  AN2 U5236 ( .A(U37_DATA4_53), .B(n9191), .Z(n9284) );
  AN2 U5237 ( .A(U37_DATA6_53), .B(n9192), .Z(n9283) );
  AN2 U5238 ( .A(U37_DATA1_53), .B(n9193), .Z(n9281) );
  OR2 U5239 ( .A(n9285), .B(n9286), .Z(n9279) );
  OR2 U5240 ( .A(n9287), .B(n9288), .Z(n9286) );
  AN2 U5241 ( .A(test_pat_seed_a[53]), .B(n9198), .Z(n9288) );
  AN2 U5242 ( .A(n9289), .B(n9199), .Z(n9287) );
  AN2 U5243 ( .A(test_pat_seed_b[53]), .B(n9201), .Z(n9285) );
  OR2 U5244 ( .A(n9290), .B(n9291), .Z(U35_Z_52) );
  OR2 U5245 ( .A(n9292), .B(n9293), .Z(n9291) );
  OR2 U5246 ( .A(n9294), .B(n9295), .Z(n9293) );
  AN2 U5247 ( .A(U37_DATA4_52), .B(n9191), .Z(n9295) );
  AN2 U5248 ( .A(U37_DATA6_52), .B(n9192), .Z(n9294) );
  AN2 U5249 ( .A(U37_DATA1_52), .B(n9193), .Z(n9292) );
  OR2 U5250 ( .A(n9296), .B(n9297), .Z(n9290) );
  OR2 U5251 ( .A(n9298), .B(n9299), .Z(n9297) );
  AN2 U5252 ( .A(test_pat_seed_a[52]), .B(n9198), .Z(n9299) );
  AN2 U5253 ( .A(n9300), .B(n9199), .Z(n9298) );
  AN2 U5254 ( .A(test_pat_seed_b[52]), .B(n9201), .Z(n9296) );
  OR2 U5255 ( .A(n9301), .B(n9302), .Z(U35_Z_51) );
  OR2 U5256 ( .A(n9303), .B(n9304), .Z(n9302) );
  OR2 U5257 ( .A(n9305), .B(n9306), .Z(n9304) );
  AN2 U5258 ( .A(U37_DATA4_51), .B(n9191), .Z(n9306) );
  AN2 U5259 ( .A(U37_DATA6_51), .B(n9192), .Z(n9305) );
  AN2 U5260 ( .A(U37_DATA1_51), .B(n9193), .Z(n9303) );
  OR2 U5261 ( .A(n9307), .B(n9308), .Z(n9301) );
  OR2 U5262 ( .A(n9309), .B(n9310), .Z(n9308) );
  AN2 U5263 ( .A(test_pat_seed_a[51]), .B(n9198), .Z(n9310) );
  AN2 U5264 ( .A(n9199), .B(n9311), .Z(n9309) );
  AN2 U5265 ( .A(test_pat_seed_b[51]), .B(n9201), .Z(n9307) );
  OR2 U5266 ( .A(n9312), .B(n9313), .Z(U35_Z_50) );
  OR2 U5267 ( .A(n9314), .B(n9315), .Z(n9313) );
  OR2 U5268 ( .A(n9316), .B(n9317), .Z(n9315) );
  AN2 U5269 ( .A(U37_DATA4_50), .B(n9191), .Z(n9317) );
  AN2 U5270 ( .A(U37_DATA6_50), .B(n9192), .Z(n9316) );
  AN2 U5271 ( .A(U37_DATA1_50), .B(n9193), .Z(n9314) );
  OR2 U5272 ( .A(n9318), .B(n9319), .Z(n9312) );
  OR2 U5273 ( .A(n9320), .B(n9321), .Z(n9319) );
  AN2 U5274 ( .A(test_pat_seed_a[50]), .B(n9198), .Z(n9321) );
  AN2 U5275 ( .A(n9322), .B(n9199), .Z(n9320) );
  AN2 U5276 ( .A(test_pat_seed_b[50]), .B(n9201), .Z(n9318) );
  OR2 U5277 ( .A(n9323), .B(n9324), .Z(U35_Z_5) );
  OR2 U5278 ( .A(n9325), .B(n9326), .Z(n9324) );
  OR2 U5279 ( .A(n9327), .B(n9328), .Z(n9326) );
  AN2 U5280 ( .A(U37_DATA4_5), .B(n9191), .Z(n9328) );
  AN2 U5281 ( .A(U37_DATA6_5), .B(n9192), .Z(n9327) );
  AN2 U5282 ( .A(U37_DATA1_5), .B(n9193), .Z(n9325) );
  OR2 U5283 ( .A(n9329), .B(n9330), .Z(n9323) );
  OR2 U5284 ( .A(n9331), .B(n9332), .Z(n9330) );
  AN2 U5285 ( .A(test_pat_seed_a[5]), .B(n9198), .Z(n9332) );
  AN2 U5286 ( .A(n9333), .B(n9199), .Z(n9331) );
  AN2 U5287 ( .A(test_pat_seed_b[5]), .B(n9201), .Z(n9329) );
  OR2 U5288 ( .A(n9334), .B(n9335), .Z(U35_Z_49) );
  OR2 U5289 ( .A(n9336), .B(n9337), .Z(n9335) );
  OR2 U5290 ( .A(n9338), .B(n9339), .Z(n9337) );
  AN2 U5291 ( .A(U37_DATA4_49), .B(n9191), .Z(n9339) );
  AN2 U5292 ( .A(U37_DATA6_49), .B(n9192), .Z(n9338) );
  AN2 U5293 ( .A(U37_DATA1_49), .B(n9193), .Z(n9336) );
  OR2 U5294 ( .A(n9340), .B(n9341), .Z(n9334) );
  OR2 U5295 ( .A(n9342), .B(n9343), .Z(n9341) );
  AN2 U5296 ( .A(test_pat_seed_a[49]), .B(n9198), .Z(n9343) );
  AN2 U5297 ( .A(n9199), .B(n9344), .Z(n9342) );
  AN2 U5298 ( .A(test_pat_seed_b[49]), .B(n9201), .Z(n9340) );
  OR2 U5299 ( .A(n9345), .B(n9346), .Z(U35_Z_48) );
  OR2 U5300 ( .A(n9347), .B(n9348), .Z(n9346) );
  OR2 U5301 ( .A(n9349), .B(n9350), .Z(n9348) );
  AN2 U5302 ( .A(U37_DATA4_48), .B(n9191), .Z(n9350) );
  AN2 U5303 ( .A(U37_DATA6_48), .B(n9192), .Z(n9349) );
  AN2 U5304 ( .A(U37_DATA1_48), .B(n9193), .Z(n9347) );
  OR2 U5305 ( .A(n9351), .B(n9352), .Z(n9345) );
  OR2 U5306 ( .A(n9353), .B(n9354), .Z(n9352) );
  AN2 U5307 ( .A(test_pat_seed_a[48]), .B(n9198), .Z(n9354) );
  AN2 U5308 ( .A(n9199), .B(n9355), .Z(n9353) );
  AN2 U5309 ( .A(test_pat_seed_b[48]), .B(n9201), .Z(n9351) );
  OR2 U5310 ( .A(n9356), .B(n9357), .Z(U35_Z_47) );
  OR2 U5311 ( .A(n9358), .B(n9359), .Z(n9357) );
  OR2 U5312 ( .A(n9360), .B(n9361), .Z(n9359) );
  AN2 U5313 ( .A(U37_DATA4_47), .B(n9191), .Z(n9361) );
  AN2 U5314 ( .A(U37_DATA6_47), .B(n9192), .Z(n9360) );
  AN2 U5315 ( .A(U37_DATA1_47), .B(n9193), .Z(n9358) );
  OR2 U5316 ( .A(n9362), .B(n9363), .Z(n9356) );
  OR2 U5317 ( .A(n9364), .B(n9365), .Z(n9363) );
  AN2 U5318 ( .A(test_pat_seed_a[47]), .B(n9198), .Z(n9365) );
  AN2 U5319 ( .A(n9199), .B(n9366), .Z(n9364) );
  AN2 U5320 ( .A(test_pat_seed_b[47]), .B(n9201), .Z(n9362) );
  OR2 U5321 ( .A(n9367), .B(n9368), .Z(U35_Z_46) );
  OR2 U5322 ( .A(n9369), .B(n9370), .Z(n9368) );
  OR2 U5323 ( .A(n9371), .B(n9372), .Z(n9370) );
  AN2 U5324 ( .A(U37_DATA4_46), .B(n9191), .Z(n9372) );
  AN2 U5325 ( .A(U37_DATA6_46), .B(n9192), .Z(n9371) );
  AN2 U5326 ( .A(U37_DATA1_46), .B(n9193), .Z(n9369) );
  OR2 U5327 ( .A(n9373), .B(n9374), .Z(n9367) );
  OR2 U5328 ( .A(n9375), .B(n9376), .Z(n9374) );
  AN2 U5329 ( .A(test_pat_seed_a[46]), .B(n9198), .Z(n9376) );
  AN2 U5330 ( .A(n9199), .B(n9377), .Z(n9375) );
  AN2 U5331 ( .A(test_pat_seed_b[46]), .B(n9201), .Z(n9373) );
  OR2 U5332 ( .A(n9378), .B(n9379), .Z(U35_Z_45) );
  OR2 U5333 ( .A(n9380), .B(n9381), .Z(n9379) );
  OR2 U5334 ( .A(n9382), .B(n9383), .Z(n9381) );
  AN2 U5335 ( .A(U37_DATA4_45), .B(n9191), .Z(n9383) );
  AN2 U5336 ( .A(U37_DATA6_45), .B(n9192), .Z(n9382) );
  AN2 U5337 ( .A(U37_DATA1_45), .B(n9193), .Z(n9380) );
  OR2 U5338 ( .A(n9384), .B(n9385), .Z(n9378) );
  OR2 U5339 ( .A(n9386), .B(n9387), .Z(n9385) );
  AN2 U5340 ( .A(test_pat_seed_a[45]), .B(n9198), .Z(n9387) );
  AN2 U5341 ( .A(n9199), .B(n9388), .Z(n9386) );
  AN2 U5342 ( .A(test_pat_seed_b[45]), .B(n9201), .Z(n9384) );
  OR2 U5343 ( .A(n9389), .B(n9390), .Z(U35_Z_44) );
  OR2 U5344 ( .A(n9391), .B(n9392), .Z(n9390) );
  OR2 U5345 ( .A(n9393), .B(n9394), .Z(n9392) );
  AN2 U5346 ( .A(U37_DATA4_44), .B(n9191), .Z(n9394) );
  AN2 U5347 ( .A(U37_DATA6_44), .B(n9192), .Z(n9393) );
  AN2 U5348 ( .A(U37_DATA1_44), .B(n9193), .Z(n9391) );
  OR2 U5349 ( .A(n9395), .B(n9396), .Z(n9389) );
  OR2 U5350 ( .A(n9397), .B(n9398), .Z(n9396) );
  AN2 U5351 ( .A(test_pat_seed_a[44]), .B(n9198), .Z(n9398) );
  AN2 U5352 ( .A(n9199), .B(n9399), .Z(n9397) );
  AN2 U5353 ( .A(test_pat_seed_b[44]), .B(n9201), .Z(n9395) );
  OR2 U5354 ( .A(n9400), .B(n9401), .Z(U35_Z_43) );
  OR2 U5355 ( .A(n9402), .B(n9403), .Z(n9401) );
  OR2 U5356 ( .A(n9404), .B(n9405), .Z(n9403) );
  AN2 U5357 ( .A(U37_DATA4_43), .B(n9191), .Z(n9405) );
  AN2 U5358 ( .A(U37_DATA6_43), .B(n9192), .Z(n9404) );
  AN2 U5359 ( .A(U37_DATA1_43), .B(n9193), .Z(n9402) );
  OR2 U5360 ( .A(n9406), .B(n9407), .Z(n9400) );
  OR2 U5361 ( .A(n9408), .B(n9409), .Z(n9407) );
  AN2 U5362 ( .A(test_pat_seed_a[43]), .B(n9198), .Z(n9409) );
  AN2 U5363 ( .A(n9199), .B(n9410), .Z(n9408) );
  AN2 U5364 ( .A(test_pat_seed_b[43]), .B(n9201), .Z(n9406) );
  OR2 U5365 ( .A(n9411), .B(n9412), .Z(U35_Z_42) );
  OR2 U5366 ( .A(n9413), .B(n9414), .Z(n9412) );
  OR2 U5367 ( .A(n9415), .B(n9416), .Z(n9414) );
  AN2 U5368 ( .A(U37_DATA4_42), .B(n9191), .Z(n9416) );
  AN2 U5369 ( .A(U37_DATA6_42), .B(n9192), .Z(n9415) );
  AN2 U5370 ( .A(U37_DATA1_42), .B(n9193), .Z(n9413) );
  OR2 U5371 ( .A(n9417), .B(n9418), .Z(n9411) );
  OR2 U5372 ( .A(n9419), .B(n9420), .Z(n9418) );
  AN2 U5373 ( .A(test_pat_seed_a[42]), .B(n9198), .Z(n9420) );
  AN2 U5374 ( .A(n9199), .B(n9421), .Z(n9419) );
  AN2 U5375 ( .A(test_pat_seed_b[42]), .B(n9201), .Z(n9417) );
  OR2 U5376 ( .A(n9422), .B(n9423), .Z(U35_Z_41) );
  OR2 U5377 ( .A(n9424), .B(n9425), .Z(n9423) );
  OR2 U5378 ( .A(n9426), .B(n9427), .Z(n9425) );
  AN2 U5379 ( .A(U37_DATA4_41), .B(n9191), .Z(n9427) );
  AN2 U5380 ( .A(U37_DATA6_41), .B(n9192), .Z(n9426) );
  AN2 U5381 ( .A(U37_DATA1_41), .B(n9193), .Z(n9424) );
  OR2 U5382 ( .A(n9428), .B(n9429), .Z(n9422) );
  OR2 U5383 ( .A(n9430), .B(n9431), .Z(n9429) );
  AN2 U5384 ( .A(test_pat_seed_a[41]), .B(n9198), .Z(n9431) );
  AN2 U5385 ( .A(n9199), .B(n9432), .Z(n9430) );
  AN2 U5386 ( .A(test_pat_seed_b[41]), .B(n9201), .Z(n9428) );
  OR2 U5387 ( .A(n9433), .B(n9434), .Z(U35_Z_40) );
  OR2 U5388 ( .A(n9435), .B(n9436), .Z(n9434) );
  OR2 U5389 ( .A(n9437), .B(n9438), .Z(n9436) );
  AN2 U5390 ( .A(U37_DATA4_40), .B(n9191), .Z(n9438) );
  AN2 U5391 ( .A(U37_DATA6_40), .B(n9192), .Z(n9437) );
  AN2 U5392 ( .A(U37_DATA1_40), .B(n9193), .Z(n9435) );
  OR2 U5393 ( .A(n9439), .B(n9440), .Z(n9433) );
  OR2 U5394 ( .A(n9441), .B(n9442), .Z(n9440) );
  AN2 U5395 ( .A(test_pat_seed_a[40]), .B(n9198), .Z(n9442) );
  AN2 U5396 ( .A(n9199), .B(n9443), .Z(n9441) );
  AN2 U5397 ( .A(test_pat_seed_b[40]), .B(n9201), .Z(n9439) );
  OR2 U5398 ( .A(n9444), .B(n9445), .Z(U35_Z_4) );
  OR2 U5399 ( .A(n9446), .B(n9447), .Z(n9445) );
  OR2 U5400 ( .A(n9448), .B(n9449), .Z(n9447) );
  AN2 U5401 ( .A(U37_DATA4_4), .B(n9191), .Z(n9449) );
  AN2 U5402 ( .A(U37_DATA6_4), .B(n9192), .Z(n9448) );
  AN2 U5403 ( .A(U37_DATA1_4), .B(n9193), .Z(n9446) );
  OR2 U5404 ( .A(n9450), .B(n9451), .Z(n9444) );
  OR2 U5405 ( .A(n9452), .B(n9453), .Z(n9451) );
  AN2 U5406 ( .A(test_pat_seed_a[4]), .B(n9198), .Z(n9453) );
  AN2 U5407 ( .A(n9199), .B(n9454), .Z(n9452) );
  AN2 U5408 ( .A(test_pat_seed_b[4]), .B(n9201), .Z(n9450) );
  OR2 U5409 ( .A(n9455), .B(n9456), .Z(U35_Z_39) );
  OR2 U5410 ( .A(n9457), .B(n9458), .Z(n9456) );
  OR2 U5411 ( .A(n9459), .B(n9460), .Z(n9458) );
  AN2 U5412 ( .A(U37_DATA4_39), .B(n9191), .Z(n9460) );
  AN2 U5413 ( .A(U37_DATA6_39), .B(n9192), .Z(n9459) );
  AN2 U5414 ( .A(U37_DATA1_39), .B(n9193), .Z(n9457) );
  OR2 U5415 ( .A(n9461), .B(n9462), .Z(n9455) );
  OR2 U5416 ( .A(n9463), .B(n9464), .Z(n9462) );
  AN2 U5417 ( .A(test_pat_seed_a[39]), .B(n9198), .Z(n9464) );
  AN2 U5418 ( .A(n9199), .B(n9465), .Z(n9463) );
  AN2 U5419 ( .A(test_pat_seed_b[39]), .B(n9201), .Z(n9461) );
  OR2 U5420 ( .A(n9466), .B(n9467), .Z(U35_Z_38) );
  OR2 U5421 ( .A(n9468), .B(n9469), .Z(n9467) );
  OR2 U5422 ( .A(n9470), .B(n9471), .Z(n9469) );
  AN2 U5423 ( .A(U37_DATA4_38), .B(n9191), .Z(n9471) );
  AN2 U5424 ( .A(U37_DATA6_38), .B(n9192), .Z(n9470) );
  AN2 U5425 ( .A(U37_DATA1_38), .B(n9193), .Z(n9468) );
  OR2 U5426 ( .A(n9472), .B(n9473), .Z(n9466) );
  OR2 U5427 ( .A(n9474), .B(n9475), .Z(n9473) );
  AN2 U5428 ( .A(test_pat_seed_a[38]), .B(n9198), .Z(n9475) );
  AN2 U5429 ( .A(n9199), .B(n9476), .Z(n9474) );
  AN2 U5430 ( .A(test_pat_seed_b[38]), .B(n9201), .Z(n9472) );
  OR2 U5431 ( .A(n9477), .B(n9478), .Z(U35_Z_37) );
  OR2 U5432 ( .A(n9479), .B(n9480), .Z(n9478) );
  OR2 U5433 ( .A(n9481), .B(n9482), .Z(n9480) );
  AN2 U5434 ( .A(U37_DATA4_37), .B(n9191), .Z(n9482) );
  AN2 U5435 ( .A(U37_DATA6_37), .B(n9192), .Z(n9481) );
  AN2 U5436 ( .A(U37_DATA1_37), .B(n9193), .Z(n9479) );
  OR2 U5437 ( .A(n9483), .B(n9484), .Z(n9477) );
  OR2 U5438 ( .A(n9485), .B(n9486), .Z(n9484) );
  AN2 U5439 ( .A(test_pat_seed_a[37]), .B(n9198), .Z(n9486) );
  AN2 U5440 ( .A(n9199), .B(n9487), .Z(n9485) );
  AN2 U5441 ( .A(test_pat_seed_b[37]), .B(n9201), .Z(n9483) );
  OR2 U5442 ( .A(n9488), .B(n9489), .Z(U35_Z_36) );
  OR2 U5443 ( .A(n9490), .B(n9491), .Z(n9489) );
  OR2 U5444 ( .A(n9492), .B(n9493), .Z(n9491) );
  AN2 U5445 ( .A(U37_DATA4_36), .B(n9191), .Z(n9493) );
  AN2 U5446 ( .A(U37_DATA6_36), .B(n9192), .Z(n9492) );
  AN2 U5447 ( .A(U37_DATA1_36), .B(n9193), .Z(n9490) );
  OR2 U5448 ( .A(n9494), .B(n9495), .Z(n9488) );
  OR2 U5449 ( .A(n9496), .B(n9497), .Z(n9495) );
  AN2 U5450 ( .A(test_pat_seed_a[36]), .B(n9198), .Z(n9497) );
  AN2 U5451 ( .A(n9199), .B(n9498), .Z(n9496) );
  AN2 U5452 ( .A(test_pat_seed_b[36]), .B(n9201), .Z(n9494) );
  OR2 U5453 ( .A(n9499), .B(n9500), .Z(U35_Z_35) );
  OR2 U5454 ( .A(n9501), .B(n9502), .Z(n9500) );
  OR2 U5455 ( .A(n9503), .B(n9504), .Z(n9502) );
  AN2 U5456 ( .A(U37_DATA4_35), .B(n9191), .Z(n9504) );
  AN2 U5457 ( .A(U37_DATA6_35), .B(n9192), .Z(n9503) );
  AN2 U5458 ( .A(U37_DATA1_35), .B(n9193), .Z(n9501) );
  OR2 U5459 ( .A(n9505), .B(n9506), .Z(n9499) );
  OR2 U5460 ( .A(n9507), .B(n9508), .Z(n9506) );
  AN2 U5461 ( .A(test_pat_seed_a[35]), .B(n9198), .Z(n9508) );
  AN2 U5462 ( .A(n9199), .B(n9509), .Z(n9507) );
  AN2 U5463 ( .A(test_pat_seed_b[35]), .B(n9201), .Z(n9505) );
  OR2 U5464 ( .A(n9510), .B(n9511), .Z(U35_Z_34) );
  OR2 U5465 ( .A(n9512), .B(n9513), .Z(n9511) );
  OR2 U5466 ( .A(n9514), .B(n9515), .Z(n9513) );
  AN2 U5467 ( .A(U37_DATA4_34), .B(n9191), .Z(n9515) );
  AN2 U5468 ( .A(U37_DATA6_34), .B(n9192), .Z(n9514) );
  AN2 U5469 ( .A(n9193), .B(U37_DATA1_34), .Z(n9512) );
  OR2 U5470 ( .A(n9516), .B(n9517), .Z(n9510) );
  OR2 U5471 ( .A(n9518), .B(n9519), .Z(n9517) );
  AN2 U5472 ( .A(test_pat_seed_a[34]), .B(n9198), .Z(n9519) );
  AN2 U5473 ( .A(n9199), .B(n9520), .Z(n9518) );
  AN2 U5474 ( .A(test_pat_seed_b[34]), .B(n9201), .Z(n9516) );
  OR2 U5475 ( .A(n9521), .B(n9522), .Z(U35_Z_33) );
  OR2 U5476 ( .A(n9523), .B(n9524), .Z(n9522) );
  OR2 U5477 ( .A(n9525), .B(n9526), .Z(n9524) );
  AN2 U5478 ( .A(U37_DATA4_33), .B(n9191), .Z(n9526) );
  AN2 U5479 ( .A(U37_DATA6_33), .B(n9192), .Z(n9525) );
  AN2 U5480 ( .A(U37_DATA1_33), .B(n9193), .Z(n9523) );
  OR2 U5481 ( .A(n9527), .B(n9528), .Z(n9521) );
  OR2 U5482 ( .A(n9529), .B(n9530), .Z(n9528) );
  AN2 U5483 ( .A(test_pat_seed_a[33]), .B(n9198), .Z(n9530) );
  AN2 U5484 ( .A(n9199), .B(n9531), .Z(n9529) );
  AN2 U5485 ( .A(test_pat_seed_b[33]), .B(n9201), .Z(n9527) );
  OR2 U5486 ( .A(n9532), .B(n9533), .Z(U35_Z_32) );
  OR2 U5487 ( .A(n9534), .B(n9535), .Z(n9533) );
  OR2 U5488 ( .A(n9536), .B(n9537), .Z(n9535) );
  AN2 U5489 ( .A(U37_DATA4_32), .B(n9191), .Z(n9537) );
  AN2 U5490 ( .A(U37_DATA6_32), .B(n9192), .Z(n9536) );
  AN2 U5491 ( .A(U37_DATA1_32), .B(n9193), .Z(n9534) );
  OR2 U5492 ( .A(n9538), .B(n9539), .Z(n9532) );
  OR2 U5493 ( .A(n9540), .B(n9541), .Z(n9539) );
  AN2 U5494 ( .A(test_pat_seed_a[32]), .B(n9198), .Z(n9541) );
  AN2 U5495 ( .A(n9199), .B(n9542), .Z(n9540) );
  AN2 U5496 ( .A(test_pat_seed_b[32]), .B(n9201), .Z(n9538) );
  OR2 U5497 ( .A(n9543), .B(n9544), .Z(U35_Z_31) );
  OR2 U5498 ( .A(n9545), .B(n9546), .Z(n9544) );
  OR2 U5499 ( .A(n9547), .B(n9548), .Z(n9546) );
  AN2 U5500 ( .A(U37_DATA4_31), .B(n9191), .Z(n9548) );
  AN2 U5501 ( .A(U37_DATA6_31), .B(n9192), .Z(n9547) );
  AN2 U5502 ( .A(U37_DATA1_31), .B(n9193), .Z(n9545) );
  OR2 U5503 ( .A(n9549), .B(n9550), .Z(n9543) );
  OR2 U5504 ( .A(n9551), .B(n9552), .Z(n9550) );
  AN2 U5505 ( .A(test_pat_seed_a[31]), .B(n9198), .Z(n9552) );
  AN2 U5506 ( .A(n9199), .B(n9553), .Z(n9551) );
  AN2 U5507 ( .A(test_pat_seed_b[31]), .B(n9201), .Z(n9549) );
  OR2 U5508 ( .A(n9554), .B(n9555), .Z(U35_Z_30) );
  OR2 U5509 ( .A(n9556), .B(n9557), .Z(n9555) );
  OR2 U5510 ( .A(n9558), .B(n9559), .Z(n9557) );
  AN2 U5511 ( .A(U37_DATA4_30), .B(n9191), .Z(n9559) );
  AN2 U5512 ( .A(U37_DATA6_30), .B(n9192), .Z(n9558) );
  AN2 U5513 ( .A(U37_DATA1_30), .B(n9193), .Z(n9556) );
  OR2 U5514 ( .A(n9560), .B(n9561), .Z(n9554) );
  OR2 U5515 ( .A(n9562), .B(n9563), .Z(n9561) );
  AN2 U5516 ( .A(test_pat_seed_a[30]), .B(n9198), .Z(n9563) );
  AN2 U5517 ( .A(n9199), .B(n9564), .Z(n9562) );
  AN2 U5518 ( .A(test_pat_seed_b[30]), .B(n9201), .Z(n9560) );
  OR2 U5519 ( .A(n9565), .B(n9566), .Z(U35_Z_3) );
  OR2 U5520 ( .A(n9567), .B(n9568), .Z(n9566) );
  OR2 U5521 ( .A(n9569), .B(n9570), .Z(n9568) );
  AN2 U5522 ( .A(U37_DATA4_3), .B(n9191), .Z(n9570) );
  AN2 U5523 ( .A(U37_DATA6_3), .B(n9192), .Z(n9569) );
  AN2 U5524 ( .A(U37_DATA1_3), .B(n9193), .Z(n9567) );
  OR2 U5525 ( .A(n9571), .B(n9572), .Z(n9565) );
  OR2 U5526 ( .A(n9573), .B(n9574), .Z(n9572) );
  AN2 U5527 ( .A(test_pat_seed_a[3]), .B(n9198), .Z(n9574) );
  AN2 U5528 ( .A(n9199), .B(n9575), .Z(n9573) );
  AN2 U5529 ( .A(test_pat_seed_b[3]), .B(n9201), .Z(n9571) );
  OR2 U5530 ( .A(n9576), .B(n9577), .Z(U35_Z_29) );
  OR2 U5531 ( .A(n9578), .B(n9579), .Z(n9577) );
  OR2 U5532 ( .A(n9580), .B(n9581), .Z(n9579) );
  AN2 U5533 ( .A(U37_DATA4_29), .B(n9191), .Z(n9581) );
  AN2 U5534 ( .A(U37_DATA6_29), .B(n9192), .Z(n9580) );
  AN2 U5535 ( .A(U37_DATA1_29), .B(n9193), .Z(n9578) );
  OR2 U5536 ( .A(n9582), .B(n9583), .Z(n9576) );
  OR2 U5537 ( .A(n9584), .B(n9585), .Z(n9583) );
  AN2 U5538 ( .A(test_pat_seed_a[29]), .B(n9198), .Z(n9585) );
  AN2 U5539 ( .A(n9199), .B(n9586), .Z(n9584) );
  AN2 U5540 ( .A(test_pat_seed_b[29]), .B(n9201), .Z(n9582) );
  OR2 U5541 ( .A(n9587), .B(n9588), .Z(U35_Z_28) );
  OR2 U5542 ( .A(n9589), .B(n9590), .Z(n9588) );
  OR2 U5543 ( .A(n9591), .B(n9592), .Z(n9590) );
  AN2 U5544 ( .A(U37_DATA4_28), .B(n9191), .Z(n9592) );
  AN2 U5545 ( .A(U37_DATA6_28), .B(n9192), .Z(n9591) );
  AN2 U5546 ( .A(U37_DATA1_28), .B(n9193), .Z(n9589) );
  OR2 U5547 ( .A(n9593), .B(n9594), .Z(n9587) );
  OR2 U5548 ( .A(n9595), .B(n9596), .Z(n9594) );
  AN2 U5549 ( .A(test_pat_seed_a[28]), .B(n9198), .Z(n9596) );
  AN2 U5550 ( .A(n9199), .B(n9597), .Z(n9595) );
  AN2 U5551 ( .A(test_pat_seed_b[28]), .B(n9201), .Z(n9593) );
  OR2 U5552 ( .A(n9598), .B(n9599), .Z(U35_Z_27) );
  OR2 U5553 ( .A(n9600), .B(n9601), .Z(n9599) );
  OR2 U5554 ( .A(n9602), .B(n9603), .Z(n9601) );
  AN2 U5555 ( .A(U37_DATA4_27), .B(n9191), .Z(n9603) );
  AN2 U5556 ( .A(U37_DATA6_27), .B(n9192), .Z(n9602) );
  AN2 U5557 ( .A(U37_DATA1_27), .B(n9193), .Z(n9600) );
  OR2 U5558 ( .A(n9604), .B(n9605), .Z(n9598) );
  OR2 U5559 ( .A(n9606), .B(n9607), .Z(n9605) );
  AN2 U5560 ( .A(test_pat_seed_a[27]), .B(n9198), .Z(n9607) );
  AN2 U5561 ( .A(n9608), .B(n9199), .Z(n9606) );
  AN2 U5562 ( .A(test_pat_seed_b[27]), .B(n9201), .Z(n9604) );
  OR2 U5563 ( .A(n9609), .B(n9610), .Z(U35_Z_26) );
  OR2 U5564 ( .A(n9611), .B(n9612), .Z(n9610) );
  OR2 U5565 ( .A(n9613), .B(n9614), .Z(n9612) );
  AN2 U5566 ( .A(U37_DATA4_26), .B(n9191), .Z(n9614) );
  AN2 U5567 ( .A(U37_DATA6_26), .B(n9192), .Z(n9613) );
  AN2 U5568 ( .A(U37_DATA1_26), .B(n9193), .Z(n9611) );
  OR2 U5569 ( .A(n9615), .B(n9616), .Z(n9609) );
  OR2 U5570 ( .A(n9617), .B(n9618), .Z(n9616) );
  AN2 U5571 ( .A(test_pat_seed_a[26]), .B(n9198), .Z(n9618) );
  AN2 U5572 ( .A(n9619), .B(n9199), .Z(n9617) );
  AN2 U5573 ( .A(test_pat_seed_b[26]), .B(n9201), .Z(n9615) );
  OR2 U5574 ( .A(n9620), .B(n9621), .Z(U35_Z_25) );
  OR2 U5575 ( .A(n9622), .B(n9623), .Z(n9621) );
  OR2 U5576 ( .A(n9624), .B(n9625), .Z(n9623) );
  AN2 U5577 ( .A(U37_DATA4_25), .B(n9191), .Z(n9625) );
  AN2 U5578 ( .A(U37_DATA6_25), .B(n9192), .Z(n9624) );
  AN2 U5579 ( .A(U37_DATA1_25), .B(n9193), .Z(n9622) );
  OR2 U5580 ( .A(n9626), .B(n9627), .Z(n9620) );
  OR2 U5581 ( .A(n9628), .B(n9629), .Z(n9627) );
  AN2 U5582 ( .A(test_pat_seed_a[25]), .B(n9198), .Z(n9629) );
  AN2 U5583 ( .A(n9199), .B(n9630), .Z(n9628) );
  AN2 U5584 ( .A(test_pat_seed_b[25]), .B(n9201), .Z(n9626) );
  OR2 U5585 ( .A(n9631), .B(n9632), .Z(U35_Z_24) );
  OR2 U5586 ( .A(n9633), .B(n9634), .Z(n9632) );
  OR2 U5587 ( .A(n9635), .B(n9636), .Z(n9634) );
  AN2 U5588 ( .A(U37_DATA4_24), .B(n9191), .Z(n9636) );
  AN2 U5589 ( .A(U37_DATA6_24), .B(n9192), .Z(n9635) );
  AN2 U5590 ( .A(U37_DATA1_24), .B(n9193), .Z(n9633) );
  OR2 U5591 ( .A(n9637), .B(n9638), .Z(n9631) );
  OR2 U5592 ( .A(n9639), .B(n9640), .Z(n9638) );
  AN2 U5593 ( .A(test_pat_seed_a[24]), .B(n9198), .Z(n9640) );
  AN2 U5594 ( .A(n9199), .B(n9641), .Z(n9639) );
  AN2 U5595 ( .A(test_pat_seed_b[24]), .B(n9201), .Z(n9637) );
  OR2 U5596 ( .A(n9642), .B(n9643), .Z(U35_Z_23) );
  OR2 U5597 ( .A(n9644), .B(n9645), .Z(n9643) );
  OR2 U5598 ( .A(n9646), .B(n9647), .Z(n9645) );
  AN2 U5599 ( .A(U37_DATA4_23), .B(n9191), .Z(n9647) );
  AN2 U5600 ( .A(U37_DATA6_23), .B(n9192), .Z(n9646) );
  AN2 U5601 ( .A(U37_DATA1_23), .B(n9193), .Z(n9644) );
  OR2 U5602 ( .A(n9648), .B(n9649), .Z(n9642) );
  OR2 U5603 ( .A(n9650), .B(n9651), .Z(n9649) );
  AN2 U5604 ( .A(test_pat_seed_a[23]), .B(n9198), .Z(n9651) );
  AN2 U5605 ( .A(n9199), .B(n9652), .Z(n9650) );
  AN2 U5606 ( .A(test_pat_seed_b[23]), .B(n9201), .Z(n9648) );
  OR2 U5607 ( .A(n9653), .B(n9654), .Z(U35_Z_22) );
  OR2 U5608 ( .A(n9655), .B(n9656), .Z(n9654) );
  OR2 U5609 ( .A(n9657), .B(n9658), .Z(n9656) );
  AN2 U5610 ( .A(U37_DATA4_22), .B(n9191), .Z(n9658) );
  AN2 U5611 ( .A(U37_DATA6_22), .B(n9192), .Z(n9657) );
  AN2 U5612 ( .A(U37_DATA1_22), .B(n9193), .Z(n9655) );
  OR2 U5613 ( .A(n9659), .B(n9660), .Z(n9653) );
  OR2 U5614 ( .A(n9661), .B(n9662), .Z(n9660) );
  AN2 U5615 ( .A(test_pat_seed_a[22]), .B(n9198), .Z(n9662) );
  AN2 U5616 ( .A(n9199), .B(n9663), .Z(n9661) );
  AN2 U5617 ( .A(test_pat_seed_b[22]), .B(n9201), .Z(n9659) );
  OR2 U5618 ( .A(n9664), .B(n9665), .Z(U35_Z_21) );
  OR2 U5619 ( .A(n9666), .B(n9667), .Z(n9665) );
  OR2 U5620 ( .A(n9668), .B(n9669), .Z(n9667) );
  AN2 U5621 ( .A(U37_DATA4_21), .B(n9191), .Z(n9669) );
  AN2 U5622 ( .A(U37_DATA6_21), .B(n9192), .Z(n9668) );
  AN2 U5623 ( .A(U37_DATA1_21), .B(n9193), .Z(n9666) );
  OR2 U5624 ( .A(n9670), .B(n9671), .Z(n9664) );
  OR2 U5625 ( .A(n9672), .B(n9673), .Z(n9671) );
  AN2 U5626 ( .A(test_pat_seed_a[21]), .B(n9198), .Z(n9673) );
  AN2 U5627 ( .A(n9199), .B(n9674), .Z(n9672) );
  AN2 U5628 ( .A(test_pat_seed_b[21]), .B(n9201), .Z(n9670) );
  OR2 U5629 ( .A(n9675), .B(n9676), .Z(U35_Z_20) );
  OR2 U5630 ( .A(n9677), .B(n9678), .Z(n9676) );
  OR2 U5631 ( .A(n9679), .B(n9680), .Z(n9678) );
  AN2 U5632 ( .A(U37_DATA4_20), .B(n9191), .Z(n9680) );
  AN2 U5633 ( .A(U37_DATA6_20), .B(n9192), .Z(n9679) );
  AN2 U5634 ( .A(U37_DATA1_20), .B(n9193), .Z(n9677) );
  OR2 U5635 ( .A(n9681), .B(n9682), .Z(n9675) );
  OR2 U5636 ( .A(n9683), .B(n9684), .Z(n9682) );
  AN2 U5637 ( .A(test_pat_seed_a[20]), .B(n9198), .Z(n9684) );
  AN2 U5638 ( .A(n9685), .B(n9199), .Z(n9683) );
  AN2 U5639 ( .A(test_pat_seed_b[20]), .B(n9201), .Z(n9681) );
  OR2 U5640 ( .A(n9686), .B(n9687), .Z(U35_Z_2) );
  OR2 U5641 ( .A(n9688), .B(n9689), .Z(n9687) );
  OR2 U5642 ( .A(n9690), .B(n9691), .Z(n9689) );
  AN2 U5643 ( .A(U37_DATA4_2), .B(n9191), .Z(n9691) );
  AN2 U5644 ( .A(U37_DATA6_2), .B(n9192), .Z(n9690) );
  AN2 U5645 ( .A(U37_DATA1_2), .B(n9193), .Z(n9688) );
  OR2 U5646 ( .A(n9692), .B(n9693), .Z(n9686) );
  OR2 U5647 ( .A(n9694), .B(n9695), .Z(n9693) );
  AN2 U5648 ( .A(test_pat_seed_a[2]), .B(n9198), .Z(n9695) );
  AN2 U5649 ( .A(n9199), .B(n9696), .Z(n9694) );
  AN2 U5650 ( .A(test_pat_seed_b[2]), .B(n9201), .Z(n9692) );
  OR2 U5651 ( .A(n9697), .B(n9698), .Z(U35_Z_19) );
  OR2 U5652 ( .A(n9699), .B(n9700), .Z(n9698) );
  OR2 U5653 ( .A(n9701), .B(n9702), .Z(n9700) );
  AN2 U5654 ( .A(U37_DATA4_19), .B(n9191), .Z(n9702) );
  AN2 U5655 ( .A(U37_DATA6_19), .B(n9192), .Z(n9701) );
  AN2 U5656 ( .A(U37_DATA1_19), .B(n9193), .Z(n9699) );
  OR2 U5657 ( .A(n9703), .B(n9704), .Z(n9697) );
  OR2 U5658 ( .A(n9705), .B(n9706), .Z(n9704) );
  AN2 U5659 ( .A(test_pat_seed_a[19]), .B(n9198), .Z(n9706) );
  AN2 U5660 ( .A(n9707), .B(n9199), .Z(n9705) );
  AN2 U5661 ( .A(test_pat_seed_b[19]), .B(n9201), .Z(n9703) );
  OR2 U5662 ( .A(n9708), .B(n9709), .Z(U35_Z_18) );
  OR2 U5663 ( .A(n9710), .B(n9711), .Z(n9709) );
  OR2 U5664 ( .A(n9712), .B(n9713), .Z(n9711) );
  AN2 U5665 ( .A(U37_DATA4_18), .B(n9191), .Z(n9713) );
  AN2 U5666 ( .A(U37_DATA6_18), .B(n9192), .Z(n9712) );
  AN2 U5667 ( .A(U37_DATA1_18), .B(n9193), .Z(n9710) );
  OR2 U5668 ( .A(n9714), .B(n9715), .Z(n9708) );
  OR2 U5669 ( .A(n9716), .B(n9717), .Z(n9715) );
  AN2 U5670 ( .A(test_pat_seed_a[18]), .B(n9198), .Z(n9717) );
  AN2 U5671 ( .A(n9718), .B(n9199), .Z(n9716) );
  AN2 U5672 ( .A(test_pat_seed_b[18]), .B(n9201), .Z(n9714) );
  OR2 U5673 ( .A(n9719), .B(n9720), .Z(U35_Z_17) );
  OR2 U5674 ( .A(n9721), .B(n9722), .Z(n9720) );
  OR2 U5675 ( .A(n9723), .B(n9724), .Z(n9722) );
  AN2 U5676 ( .A(U37_DATA4_17), .B(n9191), .Z(n9724) );
  AN2 U5677 ( .A(U37_DATA6_17), .B(n9192), .Z(n9723) );
  AN2 U5678 ( .A(U37_DATA1_17), .B(n9193), .Z(n9721) );
  OR2 U5679 ( .A(n9725), .B(n9726), .Z(n9719) );
  OR2 U5680 ( .A(n9727), .B(n9728), .Z(n9726) );
  AN2 U5681 ( .A(test_pat_seed_a[17]), .B(n9198), .Z(n9728) );
  AN2 U5682 ( .A(n9199), .B(n9729), .Z(n9727) );
  AN2 U5683 ( .A(test_pat_seed_b[17]), .B(n9201), .Z(n9725) );
  OR2 U5684 ( .A(n9730), .B(n9731), .Z(U35_Z_16) );
  OR2 U5685 ( .A(n9732), .B(n9733), .Z(n9731) );
  OR2 U5686 ( .A(n9734), .B(n9735), .Z(n9733) );
  AN2 U5687 ( .A(U37_DATA4_16), .B(n9191), .Z(n9735) );
  AN2 U5688 ( .A(U37_DATA6_16), .B(n9192), .Z(n9734) );
  AN2 U5689 ( .A(U37_DATA1_16), .B(n9193), .Z(n9732) );
  OR2 U5690 ( .A(n9736), .B(n9737), .Z(n9730) );
  OR2 U5691 ( .A(n9738), .B(n9739), .Z(n9737) );
  AN2 U5692 ( .A(test_pat_seed_a[16]), .B(n9198), .Z(n9739) );
  AN2 U5693 ( .A(n9199), .B(n9740), .Z(n9738) );
  AN2 U5694 ( .A(test_pat_seed_b[16]), .B(n9201), .Z(n9736) );
  OR2 U5695 ( .A(n9741), .B(n9742), .Z(U35_Z_15) );
  OR2 U5696 ( .A(n9743), .B(n9744), .Z(n9742) );
  OR2 U5697 ( .A(n9745), .B(n9746), .Z(n9744) );
  AN2 U5698 ( .A(U37_DATA4_15), .B(n9191), .Z(n9746) );
  AN2 U5699 ( .A(U37_DATA6_15), .B(n9192), .Z(n9745) );
  AN2 U5700 ( .A(n9193), .B(U37_DATA1_15), .Z(n9743) );
  OR2 U5701 ( .A(n9747), .B(n9748), .Z(n9741) );
  OR2 U5702 ( .A(n9749), .B(n9750), .Z(n9748) );
  AN2 U5703 ( .A(test_pat_seed_a[15]), .B(n9198), .Z(n9750) );
  AN2 U5704 ( .A(n9199), .B(n9751), .Z(n9749) );
  AN2 U5705 ( .A(test_pat_seed_b[15]), .B(n9201), .Z(n9747) );
  OR2 U5706 ( .A(n9752), .B(n9753), .Z(U35_Z_14) );
  OR2 U5707 ( .A(n9754), .B(n9755), .Z(n9753) );
  OR2 U5708 ( .A(n9756), .B(n9757), .Z(n9755) );
  AN2 U5709 ( .A(U37_DATA4_14), .B(n9191), .Z(n9757) );
  AN2 U5710 ( .A(U37_DATA6_14), .B(n9192), .Z(n9756) );
  AN2 U5711 ( .A(U37_DATA1_14), .B(n9193), .Z(n9754) );
  OR2 U5712 ( .A(n9758), .B(n9759), .Z(n9752) );
  OR2 U5713 ( .A(n9760), .B(n9761), .Z(n9759) );
  AN2 U5714 ( .A(test_pat_seed_a[14]), .B(n9198), .Z(n9761) );
  AN2 U5715 ( .A(n9199), .B(n9762), .Z(n9760) );
  AN2 U5716 ( .A(test_pat_seed_b[14]), .B(n9201), .Z(n9758) );
  OR2 U5717 ( .A(n9763), .B(n9764), .Z(U35_Z_13) );
  OR2 U5718 ( .A(n9765), .B(n9766), .Z(n9764) );
  OR2 U5719 ( .A(n9767), .B(n9768), .Z(n9766) );
  AN2 U5720 ( .A(U37_DATA4_13), .B(n9191), .Z(n9768) );
  AN2 U5721 ( .A(U37_DATA6_13), .B(n9192), .Z(n9767) );
  AN2 U5722 ( .A(U37_DATA1_13), .B(n9193), .Z(n9765) );
  OR2 U5723 ( .A(n9769), .B(n9770), .Z(n9763) );
  OR2 U5724 ( .A(n9771), .B(n9772), .Z(n9770) );
  AN2 U5725 ( .A(test_pat_seed_a[13]), .B(n9198), .Z(n9772) );
  AN2 U5726 ( .A(n9773), .B(n9199), .Z(n9771) );
  AN2 U5727 ( .A(test_pat_seed_b[13]), .B(n9201), .Z(n9769) );
  OR2 U5728 ( .A(n9774), .B(n9775), .Z(U35_Z_12) );
  OR2 U5729 ( .A(n9776), .B(n9777), .Z(n9775) );
  OR2 U5730 ( .A(n9778), .B(n9779), .Z(n9777) );
  AN2 U5731 ( .A(U37_DATA4_12), .B(n9191), .Z(n9779) );
  AN2 U5732 ( .A(U37_DATA6_12), .B(n9192), .Z(n9778) );
  AN2 U5733 ( .A(U37_DATA1_12), .B(n9193), .Z(n9776) );
  OR2 U5734 ( .A(n9780), .B(n9781), .Z(n9774) );
  OR2 U5735 ( .A(n9782), .B(n9783), .Z(n9781) );
  AN2 U5736 ( .A(test_pat_seed_a[12]), .B(n9198), .Z(n9783) );
  AN2 U5737 ( .A(n9784), .B(n9199), .Z(n9782) );
  AN2 U5738 ( .A(test_pat_seed_b[12]), .B(n9201), .Z(n9780) );
  OR2 U5739 ( .A(n9785), .B(n9786), .Z(U35_Z_11) );
  OR2 U5740 ( .A(n9787), .B(n9788), .Z(n9786) );
  OR2 U5741 ( .A(n9789), .B(n9790), .Z(n9788) );
  AN2 U5742 ( .A(U37_DATA4_11), .B(n9191), .Z(n9790) );
  AN2 U5743 ( .A(U37_DATA6_11), .B(n9192), .Z(n9789) );
  AN2 U5744 ( .A(U37_DATA1_11), .B(n9193), .Z(n9787) );
  OR2 U5745 ( .A(n9791), .B(n9792), .Z(n9785) );
  OR2 U5746 ( .A(n9793), .B(n9794), .Z(n9792) );
  AN2 U5747 ( .A(test_pat_seed_a[11]), .B(n9198), .Z(n9794) );
  AN2 U5748 ( .A(n9199), .B(n9795), .Z(n9793) );
  AN2 U5749 ( .A(test_pat_seed_b[11]), .B(n9201), .Z(n9791) );
  OR2 U5750 ( .A(n9796), .B(n9797), .Z(U35_Z_10) );
  OR2 U5751 ( .A(n9798), .B(n9799), .Z(n9797) );
  OR2 U5752 ( .A(n9800), .B(n9801), .Z(n9799) );
  AN2 U5753 ( .A(U37_DATA4_10), .B(n9191), .Z(n9801) );
  AN2 U5754 ( .A(U37_DATA6_10), .B(n9192), .Z(n9800) );
  AN2 U5755 ( .A(U37_DATA1_10), .B(n9193), .Z(n9798) );
  OR2 U5756 ( .A(n9802), .B(n9803), .Z(n9796) );
  OR2 U5757 ( .A(n9804), .B(n9805), .Z(n9803) );
  AN2 U5758 ( .A(test_pat_seed_a[10]), .B(n9198), .Z(n9805) );
  AN2 U5759 ( .A(n9199), .B(n9806), .Z(n9804) );
  AN2 U5760 ( .A(test_pat_seed_b[10]), .B(n9201), .Z(n9802) );
  OR2 U5761 ( .A(n9807), .B(n9808), .Z(U35_Z_1) );
  OR2 U5762 ( .A(n9809), .B(n9810), .Z(n9808) );
  OR2 U5763 ( .A(n9811), .B(n9812), .Z(n9810) );
  AN2 U5764 ( .A(U37_DATA4_1), .B(n9191), .Z(n9812) );
  AN2 U5765 ( .A(U37_DATA6_1), .B(n9192), .Z(n9811) );
  AN2 U5766 ( .A(U37_DATA1_1), .B(n9193), .Z(n9809) );
  OR2 U5767 ( .A(n9813), .B(n9814), .Z(n9807) );
  OR2 U5768 ( .A(n9815), .B(n9816), .Z(n9814) );
  AN2 U5769 ( .A(test_pat_seed_a[1]), .B(n9198), .Z(n9816) );
  AN2 U5770 ( .A(n9817), .B(n9199), .Z(n9815) );
  AN2 U5771 ( .A(test_pat_seed_b[1]), .B(n9201), .Z(n9813) );
  OR2 U5772 ( .A(n9818), .B(n9819), .Z(U35_Z_0) );
  OR2 U5773 ( .A(n9820), .B(n9821), .Z(n9819) );
  OR2 U5774 ( .A(n9822), .B(n9823), .Z(n9821) );
  AN2 U5775 ( .A(U37_DATA4_0), .B(n9191), .Z(n9823) );
  AN2 U5776 ( .A(n9824), .B(n9825), .Z(n9191) );
  AN2 U5777 ( .A(n9826), .B(n1256), .Z(n9825) );
  IV U5778 ( .A(n1244), .Z(n9826) );
  AN2 U5779 ( .A(U37_DATA6_0), .B(n9192), .Z(n9822) );
  AN2 U5780 ( .A(n9827), .B(n9828), .Z(n9192) );
  AN2 U5781 ( .A(n1235), .B(n1148), .Z(n9828) );
  AN2 U5782 ( .A(n9829), .B(n8648), .Z(n9827) );
  IV U5783 ( .A(n1226), .Z(n9829) );
  AN2 U5784 ( .A(U37_DATA1_0), .B(n9193), .Z(n9820) );
  OR2 U5785 ( .A(n9830), .B(n9831), .Z(n9818) );
  OR2 U5786 ( .A(n9832), .B(n9833), .Z(n9831) );
  AN2 U5787 ( .A(test_pat_seed_a[0]), .B(n9198), .Z(n9833) );
  AN2 U5788 ( .A(n9834), .B(n9824), .Z(n9198) );
  IV U5789 ( .A(n1256), .Z(n9834) );
  AN2 U5790 ( .A(n9835), .B(n9199), .Z(n9832) );
  AN2 U5791 ( .A(n1148), .B(n1935), .Z(n9199) );
  AN2 U5792 ( .A(test_pat_seed_b[0]), .B(n9201), .Z(n9830) );
  AN2 U5793 ( .A(n1148), .B(n9836), .Z(n9201) );
  AN2 U5794 ( .A(n9837), .B(n8648), .Z(n9836) );
  AN2 U5795 ( .A(n9838), .B(n9839), .Z(n8648) );
  AN2 U5796 ( .A(n1256), .B(tx_fifo_pop_2), .Z(n9839) );
  AN2 U5797 ( .A(n98), .B(n1244), .Z(n9838) );
  IV U5798 ( .A(n1235), .Z(n9837) );
  OR2 U5799 ( .A(n9840), .B(n9841), .Z(U34_Z_8) );
  AN2 U5800 ( .A(n9842), .B(n5628), .Z(n9841) );
  IV U5801 ( .A(U4_DATA1_8), .Z(n5628) );
  AN2 U5802 ( .A(n9843), .B(n9844), .Z(n9842) );
  AN2 U5803 ( .A(n9824), .B(U4_DATA1_7), .Z(n9843) );
  AN2 U5804 ( .A(n9845), .B(U4_DATA1_8), .Z(n9840) );
  OR2 U5805 ( .A(n9846), .B(n9847), .Z(n9845) );
  AN2 U5806 ( .A(n9848), .B(n5627), .Z(n9846) );
  OR2 U5807 ( .A(n9849), .B(n9850), .Z(U34_Z_7) );
  AN2 U5808 ( .A(n9851), .B(n5627), .Z(n9850) );
  IV U5809 ( .A(U4_DATA1_7), .Z(n5627) );
  AN2 U5810 ( .A(n9844), .B(n9824), .Z(n9851) );
  IV U5811 ( .A(n9852), .Z(n9844) );
  AN2 U5812 ( .A(n9847), .B(U4_DATA1_7), .Z(n9849) );
  OR2 U5813 ( .A(n9853), .B(n9854), .Z(n9847) );
  AN2 U5814 ( .A(n9848), .B(n9852), .Z(n9853) );
  OR2 U5815 ( .A(n9855), .B(n9856), .Z(n9852) );
  OR2 U5816 ( .A(n9857), .B(n9858), .Z(n9856) );
  OR2 U5817 ( .A(n9859), .B(n9860), .Z(U34_Z_6) );
  AN2 U5818 ( .A(n9861), .B(n9855), .Z(n9860) );
  IV U5819 ( .A(U4_DATA1_6), .Z(n9855) );
  AN2 U5820 ( .A(n9862), .B(U4_DATA1_5), .Z(n9861) );
  AN2 U5821 ( .A(U4_DATA1_6), .B(n9863), .Z(n9859) );
  OR2 U5822 ( .A(n9864), .B(n9865), .Z(n9863) );
  AN2 U5823 ( .A(n9848), .B(n9858), .Z(n9864) );
  OR2 U5824 ( .A(n9866), .B(n9867), .Z(U34_Z_5) );
  AN2 U5825 ( .A(n9862), .B(n9858), .Z(n9867) );
  IV U5826 ( .A(U4_DATA1_5), .Z(n9858) );
  AN2 U5827 ( .A(n9868), .B(n9824), .Z(n9862) );
  IV U5828 ( .A(n9857), .Z(n9868) );
  AN2 U5829 ( .A(U4_DATA1_5), .B(n9865), .Z(n9866) );
  OR2 U5830 ( .A(n9869), .B(n9854), .Z(n9865) );
  AN2 U5831 ( .A(n9848), .B(n9857), .Z(n9869) );
  OR2 U5832 ( .A(n9870), .B(n9871), .Z(n9857) );
  OR2 U5833 ( .A(n9872), .B(n9873), .Z(n9871) );
  OR2 U5834 ( .A(n9874), .B(n9875), .Z(U34_Z_4) );
  AN2 U5835 ( .A(n9876), .B(n9870), .Z(n9875) );
  IV U5836 ( .A(U4_DATA1_4), .Z(n9870) );
  AN2 U5837 ( .A(n9877), .B(U4_DATA1_3), .Z(n9876) );
  AN2 U5838 ( .A(U4_DATA1_4), .B(n9878), .Z(n9874) );
  OR2 U5839 ( .A(n9879), .B(n9880), .Z(n9878) );
  AN2 U5840 ( .A(n9848), .B(n9873), .Z(n9879) );
  OR2 U5841 ( .A(n9881), .B(n9882), .Z(U34_Z_3) );
  AN2 U5842 ( .A(n9877), .B(n9873), .Z(n9882) );
  IV U5843 ( .A(U4_DATA1_3), .Z(n9873) );
  AN2 U5844 ( .A(n9883), .B(n9824), .Z(n9877) );
  IV U5845 ( .A(n9872), .Z(n9883) );
  AN2 U5846 ( .A(U4_DATA1_3), .B(n9880), .Z(n9881) );
  OR2 U5847 ( .A(n9884), .B(n9854), .Z(n9880) );
  AN2 U5848 ( .A(n9848), .B(n9872), .Z(n9884) );
  OR2 U5849 ( .A(n9885), .B(n9886), .Z(n9872) );
  OR2 U5850 ( .A(n9887), .B(n9888), .Z(n9886) );
  OR2 U5851 ( .A(n9889), .B(n9890), .Z(U34_Z_2) );
  AN2 U5852 ( .A(n9891), .B(n9885), .Z(n9890) );
  IV U5853 ( .A(U4_DATA1_2), .Z(n9885) );
  AN2 U5854 ( .A(n9892), .B(U4_DATA1_1), .Z(n9891) );
  AN2 U5855 ( .A(U4_DATA1_2), .B(n9893), .Z(n9889) );
  OR2 U5856 ( .A(n9894), .B(n9895), .Z(n9893) );
  AN2 U5857 ( .A(n9848), .B(n9888), .Z(n9894) );
  OR2 U5858 ( .A(n9896), .B(n9897), .Z(U34_Z_1) );
  AN2 U5859 ( .A(n9892), .B(n9888), .Z(n9897) );
  IV U5860 ( .A(U4_DATA1_1), .Z(n9888) );
  AN2 U5861 ( .A(U4_DATA1_0), .B(n9824), .Z(n9892) );
  AN2 U5862 ( .A(U4_DATA1_1), .B(n9895), .Z(n9896) );
  OR2 U5863 ( .A(n9898), .B(n9854), .Z(n9895) );
  AN2 U5864 ( .A(n98), .B(n9193), .Z(n9854) );
  AN2 U5865 ( .A(n9899), .B(n1148), .Z(n9193) );
  AN2 U5866 ( .A(n9848), .B(n9887), .Z(n9898) );
  OR2 U5867 ( .A(n9900), .B(n9901), .Z(U34_Z_0) );
  AN2 U5868 ( .A(n9902), .B(U4_DATA1_0), .Z(n9901) );
  AN2 U5869 ( .A(n9848), .B(n9899), .Z(n9902) );
  IV U5870 ( .A(tx_fifo_pop_2), .Z(n9899) );
  AN2 U5871 ( .A(n9824), .B(n9887), .Z(n9900) );
  IV U5872 ( .A(U4_DATA1_0), .Z(n9887) );
  AN2 U5873 ( .A(tx_fifo_pop_2), .B(n9848), .Z(n9824) );
  AN2 U5874 ( .A(n98), .B(n1148), .Z(n9848) );
  OR2 U5875 ( .A(n9903), .B(n9904), .Z(U3_U1_Z_9) );
  AN2 U5876 ( .A(U3_U1_DATA1_9), .B(n8661), .Z(n9904) );
  AN2 U5877 ( .A(U3_U1_DATA3_9), .B(n8662), .Z(n9903) );
  OR2 U5878 ( .A(n9905), .B(n9906), .Z(U3_U1_Z_8) );
  AN2 U5879 ( .A(U3_U1_DATA1_8), .B(n8661), .Z(n9906) );
  AN2 U5880 ( .A(U3_U1_DATA3_8), .B(n8662), .Z(n9905) );
  OR2 U5881 ( .A(n9907), .B(n9908), .Z(U3_U1_Z_7) );
  AN2 U5882 ( .A(U3_U1_DATA1_7), .B(n8661), .Z(n9908) );
  AN2 U5883 ( .A(U3_U1_DATA3_7), .B(n8662), .Z(n9907) );
  OR2 U5884 ( .A(n9909), .B(n9910), .Z(U3_U1_Z_6) );
  AN2 U5885 ( .A(U3_U1_DATA1_6), .B(n8661), .Z(n9910) );
  AN2 U5886 ( .A(U3_U1_DATA3_6), .B(n8662), .Z(n9909) );
  OR2 U5887 ( .A(n9911), .B(n9912), .Z(U3_U1_Z_5) );
  AN2 U5888 ( .A(U3_U1_DATA1_5), .B(n8661), .Z(n9912) );
  AN2 U5889 ( .A(U3_U1_DATA3_5), .B(n8662), .Z(n9911) );
  OR2 U5890 ( .A(n9913), .B(n9914), .Z(U3_U1_Z_4) );
  AN2 U5891 ( .A(U3_U1_DATA1_4), .B(n8661), .Z(n9914) );
  AN2 U5892 ( .A(U3_U1_DATA3_4), .B(n8662), .Z(n9913) );
  OR2 U5893 ( .A(n9915), .B(n9916), .Z(U3_U1_Z_3) );
  AN2 U5894 ( .A(U3_U1_DATA1_3), .B(n8661), .Z(n9916) );
  AN2 U5895 ( .A(U3_U1_DATA3_3), .B(n8662), .Z(n9915) );
  OR2 U5896 ( .A(n9917), .B(n9918), .Z(U3_U1_Z_2) );
  AN2 U5897 ( .A(U3_U1_DATA1_2), .B(n8661), .Z(n9918) );
  AN2 U5898 ( .A(U3_U1_DATA3_2), .B(n8662), .Z(n9917) );
  AN2 U5899 ( .A(U3_U1_DATA1_15), .B(n8661), .Z(U3_U1_Z_15) );
  AN2 U5900 ( .A(U3_U1_DATA1_14), .B(n8661), .Z(U3_U1_Z_14) );
  AN2 U5901 ( .A(U3_U1_DATA1_13), .B(n8661), .Z(U3_U1_Z_13) );
  AN2 U5902 ( .A(U3_U1_DATA1_12), .B(n8661), .Z(U3_U1_Z_12) );
  AN2 U5903 ( .A(U3_U1_DATA1_11), .B(n8661), .Z(U3_U1_Z_11) );
  OR2 U5904 ( .A(n9919), .B(n9920), .Z(U3_U1_Z_10) );
  AN2 U5905 ( .A(U3_U1_DATA1_10), .B(n8661), .Z(n9920) );
  AN2 U5906 ( .A(U3_U1_DATA3_10), .B(n8662), .Z(n9919) );
  OR2 U5907 ( .A(n9921), .B(n9922), .Z(U3_U1_Z_1) );
  AN2 U5908 ( .A(U3_U1_DATA1_1), .B(n8661), .Z(n9922) );
  OR2 U5909 ( .A(n9024), .B(n8719), .Z(n8661) );
  AN2 U5910 ( .A(n2549), .B(n2548), .Z(n9024) );
  AN2 U5911 ( .A(U3_U1_DATA3_1), .B(n8662), .Z(n9921) );
  IV U5912 ( .A(n9923), .Z(n8662) );
  OR2 U5913 ( .A(n2536), .B(n2537), .Z(n9923) );
  OR2 U5914 ( .A(n9924), .B(n9925), .Z(tx_data_out[9]) );
  OR2 U5915 ( .A(n9926), .B(n9927), .Z(n9925) );
  AN2 U5916 ( .A(n9928), .B(U157_Z_2), .Z(n9927) );
  AN2 U5917 ( .A(n9929), .B(n9817), .Z(n9926) );
  AN2 U5918 ( .A(n9930), .B(U40_DATA2_7), .Z(n9924) );
  OR2 U5919 ( .A(n9931), .B(n9932), .Z(tx_data_out[8]) );
  OR2 U5920 ( .A(n9933), .B(n9934), .Z(n9932) );
  AN2 U5921 ( .A(n9928), .B(U156_Z_1), .Z(n9934) );
  AN2 U5922 ( .A(n9929), .B(n9835), .Z(n9933) );
  AN2 U5923 ( .A(n9930), .B(U40_DATA2_6), .Z(n9931) );
  OR2 U5924 ( .A(n9935), .B(n9936), .Z(tx_data_out[7]) );
  OR2 U5925 ( .A(n9937), .B(n9938), .Z(n9936) );
  AN2 U5926 ( .A(n9928), .B(U156_Z_0), .Z(n9938) );
  AN2 U5927 ( .A(n9929), .B(n9939), .Z(n9937) );
  AN2 U5928 ( .A(n9930), .B(U40_DATA2_5), .Z(n9935) );
  OR2 U5929 ( .A(n9940), .B(n9941), .Z(tx_data_out[65]) );
  AN2 U5930 ( .A(n9942), .B(n9943), .Z(n9941) );
  AN2 U5931 ( .A(n9929), .B(n9245), .Z(n9940) );
  AN2 U5932 ( .A(n9944), .B(n9945), .Z(n9245) );
  OR2 U5933 ( .A(n9939), .B(n9946), .Z(n9945) );
  OR2 U5934 ( .A(n9947), .B(n9948), .Z(n9944) );
  IV U5935 ( .A(n9946), .Z(n9947) );
  OR2 U5936 ( .A(n9949), .B(n9950), .Z(n9946) );
  AN2 U5937 ( .A(n9718), .B(n9951), .Z(n9950) );
  OR2 U5938 ( .A(n9952), .B(n9953), .Z(n9951) );
  AN2 U5939 ( .A(n9954), .B(n9955), .Z(n9952) );
  IV U5940 ( .A(n9943), .Z(n9954) );
  AN2 U5941 ( .A(n9956), .B(n9957), .Z(n9949) );
  OR2 U5942 ( .A(n9958), .B(n1934), .Z(n9957) );
  AN2 U5943 ( .A(n9943), .B(n5684), .Z(n9958) );
  OR2 U5944 ( .A(n9959), .B(n9960), .Z(n9943) );
  OR2 U5945 ( .A(n9961), .B(n9962), .Z(n9960) );
  AN2 U5946 ( .A(n9963), .B(U156_Z_28), .Z(n9962) );
  AN2 U5947 ( .A(n9964), .B(n9965), .Z(n9961) );
  OR2 U5948 ( .A(n8766), .B(n9966), .Z(n9964) );
  OR2 U5949 ( .A(n8763), .B(n9967), .Z(n9966) );
  AN2 U5950 ( .A(n9968), .B(U156_Z_33), .Z(n9959) );
  OR2 U5951 ( .A(n9969), .B(n9970), .Z(tx_data_out[64]) );
  AN2 U5952 ( .A(n9942), .B(n9971), .Z(n9970) );
  AN2 U5953 ( .A(n9929), .B(n9256), .Z(n9969) );
  AN2 U5954 ( .A(n9972), .B(n9973), .Z(n9256) );
  OR2 U5955 ( .A(n9974), .B(n9975), .Z(n9973) );
  OR2 U5956 ( .A(n9976), .B(n9977), .Z(n9972) );
  IV U5957 ( .A(n9975), .Z(n9976) );
  OR2 U5958 ( .A(n9978), .B(n9979), .Z(n9975) );
  AN2 U5959 ( .A(n9729), .B(n9980), .Z(n9979) );
  OR2 U5960 ( .A(n9981), .B(n9953), .Z(n9980) );
  AN2 U5961 ( .A(n9982), .B(n9955), .Z(n9981) );
  IV U5962 ( .A(n9971), .Z(n9982) );
  AN2 U5963 ( .A(n9983), .B(n9984), .Z(n9978) );
  OR2 U5964 ( .A(n9985), .B(n1934), .Z(n9984) );
  AN2 U5965 ( .A(n9971), .B(n5684), .Z(n9985) );
  OR2 U5966 ( .A(n9986), .B(n9987), .Z(n9971) );
  OR2 U5967 ( .A(n9988), .B(n9989), .Z(n9987) );
  AN2 U5968 ( .A(n9968), .B(U156_Z_32), .Z(n9989) );
  AN2 U5969 ( .A(n9963), .B(U156_Z_27), .Z(n9988) );
  OR2 U5970 ( .A(n9990), .B(n9991), .Z(n9986) );
  AN2 U5971 ( .A(n9992), .B(n9965), .Z(n9991) );
  OR2 U5972 ( .A(n8767), .B(n9967), .Z(n9992) );
  AN2 U5973 ( .A(n9993), .B(n8770), .Z(n9967) );
  IV U5974 ( .A(n9729), .Z(n9983) );
  OR2 U5975 ( .A(n9994), .B(n9995), .Z(tx_data_out[63]) );
  AN2 U5976 ( .A(n9942), .B(n9996), .Z(n9995) );
  AN2 U5977 ( .A(n9929), .B(n9267), .Z(n9994) );
  AN2 U5978 ( .A(n9997), .B(n9998), .Z(n9267) );
  OR2 U5979 ( .A(n9999), .B(n10000), .Z(n9998) );
  OR2 U5980 ( .A(n10001), .B(n10002), .Z(n9997) );
  IV U5981 ( .A(n10000), .Z(n10001) );
  OR2 U5982 ( .A(n10003), .B(n10004), .Z(n10000) );
  AN2 U5983 ( .A(n9740), .B(n10005), .Z(n10004) );
  OR2 U5984 ( .A(n10006), .B(n9953), .Z(n10005) );
  AN2 U5985 ( .A(n10007), .B(n9955), .Z(n10006) );
  IV U5986 ( .A(n9996), .Z(n10007) );
  AN2 U5987 ( .A(n10008), .B(n10009), .Z(n10003) );
  OR2 U5988 ( .A(n10010), .B(n1934), .Z(n10009) );
  AN2 U5989 ( .A(n9996), .B(n5684), .Z(n10010) );
  OR2 U5990 ( .A(n10011), .B(n10012), .Z(n9996) );
  OR2 U5991 ( .A(n10013), .B(n10014), .Z(n10012) );
  AN2 U5992 ( .A(n9968), .B(U156_Z_31), .Z(n10013) );
  OR2 U5993 ( .A(n10015), .B(n10016), .Z(n10011) );
  AN2 U5994 ( .A(n9963), .B(U156_Z_26), .Z(n10016) );
  IV U5995 ( .A(n9740), .Z(n10008) );
  OR2 U5996 ( .A(n10017), .B(n10018), .Z(tx_data_out[62]) );
  AN2 U5997 ( .A(n9942), .B(n10019), .Z(n10018) );
  AN2 U5998 ( .A(n9929), .B(n9278), .Z(n10017) );
  AN2 U5999 ( .A(n10020), .B(n10021), .Z(n9278) );
  OR2 U6000 ( .A(n10022), .B(n10023), .Z(n10021) );
  OR2 U6001 ( .A(n10024), .B(n10025), .Z(n10020) );
  IV U6002 ( .A(n10023), .Z(n10024) );
  OR2 U6003 ( .A(n10026), .B(n10027), .Z(n10023) );
  AN2 U6004 ( .A(n9751), .B(n10028), .Z(n10027) );
  OR2 U6005 ( .A(n10029), .B(n9953), .Z(n10028) );
  AN2 U6006 ( .A(n10030), .B(n9955), .Z(n10029) );
  IV U6007 ( .A(n10019), .Z(n10030) );
  AN2 U6008 ( .A(n10031), .B(n10032), .Z(n10026) );
  OR2 U6009 ( .A(n10033), .B(n1934), .Z(n10032) );
  AN2 U6010 ( .A(n10019), .B(n5684), .Z(n10033) );
  OR2 U6011 ( .A(n10034), .B(n10035), .Z(n10019) );
  OR2 U6012 ( .A(n10014), .B(n10036), .Z(n10035) );
  OR2 U6013 ( .A(n10037), .B(n10038), .Z(n10014) );
  AN2 U6014 ( .A(n10039), .B(n9965), .Z(n10037) );
  OR2 U6015 ( .A(n10040), .B(n10041), .Z(n10039) );
  AN2 U6016 ( .A(n8721), .B(n10042), .Z(n10041) );
  OR2 U6017 ( .A(n1298), .B(n5443), .Z(n10042) );
  IV U6018 ( .A(n1397), .Z(n5443) );
  AN2 U6019 ( .A(n10043), .B(n8770), .Z(n8721) );
  IV U6020 ( .A(n9993), .Z(n10043) );
  OR2 U6021 ( .A(n5442), .B(n5436), .Z(n9993) );
  IV U6022 ( .A(n1533), .Z(n5442) );
  AN2 U6023 ( .A(n10044), .B(n8770), .Z(n10040) );
  AN2 U6024 ( .A(n1589), .B(n10045), .Z(n8770) );
  AN2 U6025 ( .A(n1533), .B(n5436), .Z(n10044) );
  IV U6026 ( .A(n1474), .Z(n5436) );
  OR2 U6027 ( .A(n10046), .B(n10047), .Z(n10034) );
  AN2 U6028 ( .A(n9968), .B(U156_Z_30), .Z(n10047) );
  AN2 U6029 ( .A(n9963), .B(U156_Z_25), .Z(n10046) );
  IV U6030 ( .A(n9751), .Z(n10031) );
  OR2 U6031 ( .A(n10048), .B(n10049), .Z(tx_data_out[61]) );
  AN2 U6032 ( .A(n9942), .B(n10050), .Z(n10049) );
  AN2 U6033 ( .A(n9929), .B(n9289), .Z(n10048) );
  AN2 U6034 ( .A(n10051), .B(n10052), .Z(n9289) );
  OR2 U6035 ( .A(n10053), .B(n10054), .Z(n10052) );
  OR2 U6036 ( .A(n10055), .B(n10056), .Z(n10051) );
  IV U6037 ( .A(n10054), .Z(n10055) );
  OR2 U6038 ( .A(n10057), .B(n10058), .Z(n10054) );
  AN2 U6039 ( .A(n9762), .B(n10059), .Z(n10058) );
  OR2 U6040 ( .A(n10060), .B(n9953), .Z(n10059) );
  AN2 U6041 ( .A(n10061), .B(n9955), .Z(n10060) );
  IV U6042 ( .A(n10050), .Z(n10061) );
  AN2 U6043 ( .A(n10062), .B(n10063), .Z(n10057) );
  OR2 U6044 ( .A(n10064), .B(n1934), .Z(n10063) );
  AN2 U6045 ( .A(n10050), .B(n5684), .Z(n10064) );
  OR2 U6046 ( .A(n10065), .B(n10066), .Z(n10050) );
  OR2 U6047 ( .A(n10067), .B(n10068), .Z(n10066) );
  AN2 U6048 ( .A(n9968), .B(U156_Z_29), .Z(n10068) );
  AN2 U6049 ( .A(n9963), .B(U156_Z_24), .Z(n10067) );
  OR2 U6050 ( .A(n10038), .B(n10069), .Z(n10065) );
  AN2 U6051 ( .A(U61_DATA2_23), .B(n9965), .Z(n10069) );
  IV U6052 ( .A(n9762), .Z(n10062) );
  OR2 U6053 ( .A(n10070), .B(n10071), .Z(tx_data_out[60]) );
  AN2 U6054 ( .A(n9942), .B(n10072), .Z(n10071) );
  AN2 U6055 ( .A(n9929), .B(n9300), .Z(n10070) );
  AN2 U6056 ( .A(n10073), .B(n10074), .Z(n9300) );
  OR2 U6057 ( .A(n10075), .B(n10076), .Z(n10074) );
  OR2 U6058 ( .A(n10077), .B(n10078), .Z(n10073) );
  IV U6059 ( .A(n10076), .Z(n10077) );
  OR2 U6060 ( .A(n10079), .B(n10080), .Z(n10076) );
  AN2 U6061 ( .A(n9773), .B(n10081), .Z(n10080) );
  OR2 U6062 ( .A(n10082), .B(n9953), .Z(n10081) );
  AN2 U6063 ( .A(n10083), .B(n9955), .Z(n10082) );
  IV U6064 ( .A(n10072), .Z(n10083) );
  AN2 U6065 ( .A(n10084), .B(n10085), .Z(n10079) );
  OR2 U6066 ( .A(n10086), .B(n1934), .Z(n10085) );
  AN2 U6067 ( .A(n10072), .B(n5684), .Z(n10086) );
  OR2 U6068 ( .A(n10087), .B(n10088), .Z(n10072) );
  OR2 U6069 ( .A(n10089), .B(n10090), .Z(n10088) );
  AN2 U6070 ( .A(n9968), .B(n8667), .Z(n10090) );
  OR2 U6071 ( .A(n4170), .B(n10091), .Z(n8667) );
  AN2 U6072 ( .A(U162_DATA3_58), .B(n10092), .Z(n10091) );
  AN2 U6073 ( .A(n9963), .B(n8668), .Z(n10089) );
  OR2 U6074 ( .A(n10038), .B(n10093), .Z(n10087) );
  AN2 U6075 ( .A(U61_DATA2_22), .B(n9965), .Z(n10093) );
  OR2 U6076 ( .A(n10094), .B(n10095), .Z(tx_data_out[6]) );
  OR2 U6077 ( .A(n10096), .B(n10097), .Z(n10095) );
  AN2 U6078 ( .A(n9928), .B(U157_Z_1), .Z(n10097) );
  AN2 U6079 ( .A(n9929), .B(n9974), .Z(n10096) );
  AN2 U6080 ( .A(n9930), .B(U40_DATA2_4), .Z(n10094) );
  OR2 U6081 ( .A(n10098), .B(n10099), .Z(tx_data_out[59]) );
  AN2 U6082 ( .A(n9942), .B(n10100), .Z(n10099) );
  AN2 U6083 ( .A(n9929), .B(n9311), .Z(n10098) );
  OR2 U6084 ( .A(n10101), .B(n10102), .Z(n9311) );
  AN2 U6085 ( .A(n10103), .B(n10104), .Z(n10102) );
  AN2 U6086 ( .A(n10105), .B(U37_DATA1_57), .Z(n10101) );
  IV U6087 ( .A(n10103), .Z(n10105) );
  OR2 U6088 ( .A(n10106), .B(n10107), .Z(n10103) );
  AN2 U6089 ( .A(n9784), .B(n10108), .Z(n10107) );
  OR2 U6090 ( .A(n10109), .B(n9953), .Z(n10108) );
  AN2 U6091 ( .A(n10110), .B(n9955), .Z(n10109) );
  IV U6092 ( .A(n10100), .Z(n10110) );
  AN2 U6093 ( .A(n10111), .B(n10112), .Z(n10106) );
  OR2 U6094 ( .A(n10113), .B(n1934), .Z(n10112) );
  AN2 U6095 ( .A(n10100), .B(n5684), .Z(n10113) );
  OR2 U6096 ( .A(n10114), .B(n10115), .Z(n10100) );
  OR2 U6097 ( .A(n10116), .B(n10036), .Z(n10115) );
  OR2 U6098 ( .A(n10117), .B(n9990), .Z(n10036) );
  AN2 U6099 ( .A(n9965), .B(n8764), .Z(n9990) );
  AN2 U6100 ( .A(n10118), .B(n10119), .Z(n8764) );
  AN2 U6101 ( .A(n5440), .B(n1696), .Z(n10119) );
  IV U6102 ( .A(n1642), .Z(n5440) );
  AN2 U6103 ( .A(n8766), .B(n9965), .Z(n10117) );
  AN2 U6104 ( .A(U154_Z_5), .B(n10120), .Z(n8766) );
  AN2 U6105 ( .A(n5438), .B(n1806), .Z(n10120) );
  IV U6106 ( .A(n1760), .Z(n5438) );
  AN2 U6107 ( .A(n9968), .B(U158_Z_14), .Z(n10116) );
  OR2 U6108 ( .A(n10015), .B(n10121), .Z(n10114) );
  AN2 U6109 ( .A(n9963), .B(U158_Z_11), .Z(n10121) );
  AN2 U6110 ( .A(n10122), .B(n9965), .Z(n10015) );
  OR2 U6111 ( .A(n10123), .B(n10124), .Z(n9965) );
  AN2 U6112 ( .A(n1930), .B(n10125), .Z(n10123) );
  OR2 U6113 ( .A(n8767), .B(n8763), .Z(n10122) );
  AN2 U6114 ( .A(n5439), .B(n10118), .Z(n8763) );
  IV U6115 ( .A(n1696), .Z(n5439) );
  AN2 U6116 ( .A(n5441), .B(n10045), .Z(n8767) );
  AN2 U6117 ( .A(n10118), .B(n10126), .Z(n10045) );
  AN2 U6118 ( .A(n1642), .B(n1696), .Z(n10126) );
  AN2 U6119 ( .A(U154_Z_5), .B(n10127), .Z(n10118) );
  AN2 U6120 ( .A(n1760), .B(n1806), .Z(n10127) );
  IV U6121 ( .A(n1589), .Z(n5441) );
  IV U6122 ( .A(n9784), .Z(n10111) );
  OR2 U6123 ( .A(n10128), .B(n10129), .Z(tx_data_out[58]) );
  AN2 U6124 ( .A(n9942), .B(n10130), .Z(n10129) );
  AN2 U6125 ( .A(n9929), .B(n9322), .Z(n10128) );
  AN2 U6126 ( .A(n10131), .B(n10132), .Z(n9322) );
  OR2 U6127 ( .A(n10133), .B(n9795), .Z(n10132) );
  IV U6128 ( .A(n10134), .Z(n10131) );
  AN2 U6129 ( .A(n9795), .B(n10133), .Z(n10134) );
  IV U6130 ( .A(n10135), .Z(n10133) );
  OR2 U6131 ( .A(n10136), .B(n10137), .Z(n10135) );
  AN2 U6132 ( .A(n10138), .B(n10139), .Z(n10137) );
  IV U6133 ( .A(n10140), .Z(n10138) );
  AN2 U6134 ( .A(U37_DATA1_56), .B(n10140), .Z(n10136) );
  OR2 U6135 ( .A(n10141), .B(n1932), .Z(n10140) );
  AN2 U6136 ( .A(n10130), .B(n5684), .Z(n10141) );
  OR2 U6137 ( .A(n10142), .B(n10143), .Z(n10130) );
  OR2 U6138 ( .A(n10144), .B(n10145), .Z(n10143) );
  AN2 U6139 ( .A(n9963), .B(U159_Z_7), .Z(n10145) );
  AN2 U6140 ( .A(n10125), .B(n5245), .Z(n9963) );
  AN2 U6141 ( .A(n10146), .B(n10147), .Z(n10144) );
  OR2 U6142 ( .A(n8777), .B(n10148), .Z(n10146) );
  OR2 U6143 ( .A(n8774), .B(n10149), .Z(n10148) );
  AN2 U6144 ( .A(n9968), .B(U158_Z_13), .Z(n10142) );
  OR2 U6145 ( .A(n10150), .B(n10151), .Z(tx_data_out[57]) );
  AN2 U6146 ( .A(n9942), .B(n10152), .Z(n10151) );
  AN2 U6147 ( .A(n9929), .B(n9344), .Z(n10150) );
  OR2 U6148 ( .A(n10153), .B(n10154), .Z(n9344) );
  AN2 U6149 ( .A(n10155), .B(n10156), .Z(n10154) );
  AN2 U6150 ( .A(n10157), .B(U37_DATA1_55), .Z(n10153) );
  IV U6151 ( .A(n10155), .Z(n10157) );
  OR2 U6152 ( .A(n10158), .B(n10159), .Z(n10155) );
  AN2 U6153 ( .A(n9806), .B(n10160), .Z(n10159) );
  OR2 U6154 ( .A(n10161), .B(n9953), .Z(n10160) );
  AN2 U6155 ( .A(n10162), .B(n9955), .Z(n10161) );
  IV U6156 ( .A(n10152), .Z(n10162) );
  AN2 U6157 ( .A(n10163), .B(n10164), .Z(n10158) );
  OR2 U6158 ( .A(n10165), .B(n1934), .Z(n10164) );
  AN2 U6159 ( .A(n10152), .B(n5684), .Z(n10165) );
  OR2 U6160 ( .A(n10166), .B(n10167), .Z(n10152) );
  OR2 U6161 ( .A(n10168), .B(n10169), .Z(n10167) );
  AN2 U6162 ( .A(n9968), .B(U156_Z_28), .Z(n10169) );
  AN2 U6163 ( .A(n10170), .B(U156_Z_23), .Z(n10168) );
  OR2 U6164 ( .A(n10171), .B(n10172), .Z(n10166) );
  AN2 U6165 ( .A(n10173), .B(n10147), .Z(n10172) );
  OR2 U6166 ( .A(n8778), .B(n10149), .Z(n10173) );
  AN2 U6167 ( .A(n10174), .B(n8781), .Z(n10149) );
  IV U6168 ( .A(n9806), .Z(n10163) );
  OR2 U6169 ( .A(n10175), .B(n10176), .Z(tx_data_out[56]) );
  AN2 U6170 ( .A(n9942), .B(n10177), .Z(n10176) );
  AN2 U6171 ( .A(n9929), .B(n9355), .Z(n10175) );
  OR2 U6172 ( .A(n10178), .B(n10179), .Z(n9355) );
  AN2 U6173 ( .A(n10180), .B(n10181), .Z(n10179) );
  AN2 U6174 ( .A(n10182), .B(U37_DATA1_54), .Z(n10178) );
  IV U6175 ( .A(n10180), .Z(n10182) );
  OR2 U6176 ( .A(n10183), .B(n10184), .Z(n10180) );
  AN2 U6177 ( .A(n9200), .B(n10185), .Z(n10184) );
  OR2 U6178 ( .A(n10186), .B(n9953), .Z(n10185) );
  AN2 U6179 ( .A(n10187), .B(n9955), .Z(n10186) );
  IV U6180 ( .A(n10177), .Z(n10187) );
  AN2 U6181 ( .A(n10188), .B(n10189), .Z(n10183) );
  OR2 U6182 ( .A(n10190), .B(n1934), .Z(n10189) );
  AN2 U6183 ( .A(n10177), .B(n5684), .Z(n10190) );
  OR2 U6184 ( .A(n10191), .B(n10192), .Z(n10177) );
  OR2 U6185 ( .A(n10193), .B(n10194), .Z(n10192) );
  AN2 U6186 ( .A(n9968), .B(U156_Z_27), .Z(n10193) );
  OR2 U6187 ( .A(n10195), .B(n10196), .Z(n10191) );
  AN2 U6188 ( .A(n10170), .B(U156_Z_22), .Z(n10196) );
  IV U6189 ( .A(n9200), .Z(n10188) );
  OR2 U6190 ( .A(n10197), .B(n10198), .Z(tx_data_out[55]) );
  AN2 U6191 ( .A(n9942), .B(n10199), .Z(n10198) );
  AN2 U6192 ( .A(n9929), .B(n9366), .Z(n10197) );
  OR2 U6193 ( .A(n10200), .B(n10201), .Z(n9366) );
  AN2 U6194 ( .A(n10202), .B(n10203), .Z(n10201) );
  AN2 U6195 ( .A(n10204), .B(U37_DATA1_53), .Z(n10200) );
  IV U6196 ( .A(n10202), .Z(n10204) );
  OR2 U6197 ( .A(n10205), .B(n10206), .Z(n10202) );
  AN2 U6198 ( .A(n9212), .B(n10207), .Z(n10206) );
  OR2 U6199 ( .A(n10208), .B(n9953), .Z(n10207) );
  AN2 U6200 ( .A(n10209), .B(n9955), .Z(n10208) );
  IV U6201 ( .A(n10199), .Z(n10209) );
  AN2 U6202 ( .A(n10210), .B(n10211), .Z(n10205) );
  OR2 U6203 ( .A(n10212), .B(n1934), .Z(n10211) );
  AN2 U6204 ( .A(n10199), .B(n5684), .Z(n10212) );
  OR2 U6205 ( .A(n10213), .B(n10214), .Z(n10199) );
  OR2 U6206 ( .A(n10194), .B(n10215), .Z(n10214) );
  OR2 U6207 ( .A(n10216), .B(n10038), .Z(n10194) );
  AN2 U6208 ( .A(n10217), .B(n10147), .Z(n10216) );
  OR2 U6209 ( .A(n10218), .B(n10219), .Z(n10217) );
  AN2 U6210 ( .A(n8723), .B(n10220), .Z(n10219) );
  OR2 U6211 ( .A(n1318), .B(n5425), .Z(n10220) );
  IV U6212 ( .A(n1423), .Z(n5425) );
  AN2 U6213 ( .A(n10221), .B(n8781), .Z(n8723) );
  IV U6214 ( .A(n10174), .Z(n10221) );
  OR2 U6215 ( .A(n5424), .B(n5418), .Z(n10174) );
  IV U6216 ( .A(n1547), .Z(n5424) );
  AN2 U6217 ( .A(n10222), .B(n8781), .Z(n10218) );
  AN2 U6218 ( .A(n1603), .B(n10223), .Z(n8781) );
  AN2 U6219 ( .A(n1547), .B(n5418), .Z(n10222) );
  IV U6220 ( .A(n1486), .Z(n5418) );
  OR2 U6221 ( .A(n10224), .B(n10225), .Z(n10213) );
  AN2 U6222 ( .A(n9968), .B(U156_Z_26), .Z(n10225) );
  AN2 U6223 ( .A(n10170), .B(U156_Z_21), .Z(n10224) );
  IV U6224 ( .A(n9212), .Z(n10210) );
  OR2 U6225 ( .A(n10226), .B(n10227), .Z(tx_data_out[54]) );
  AN2 U6226 ( .A(n9942), .B(n10228), .Z(n10227) );
  AN2 U6227 ( .A(n9929), .B(n9377), .Z(n10226) );
  OR2 U6228 ( .A(n10229), .B(n10230), .Z(n9377) );
  AN2 U6229 ( .A(n10231), .B(n10232), .Z(n10230) );
  AN2 U6230 ( .A(n10233), .B(U37_DATA1_52), .Z(n10229) );
  IV U6231 ( .A(n10231), .Z(n10233) );
  OR2 U6232 ( .A(n10234), .B(n10235), .Z(n10231) );
  AN2 U6233 ( .A(n9223), .B(n10236), .Z(n10235) );
  OR2 U6234 ( .A(n10237), .B(n9953), .Z(n10236) );
  AN2 U6235 ( .A(n10238), .B(n9955), .Z(n10237) );
  IV U6236 ( .A(n10228), .Z(n10238) );
  AN2 U6237 ( .A(n10239), .B(n10240), .Z(n10234) );
  OR2 U6238 ( .A(n10241), .B(n1934), .Z(n10240) );
  AN2 U6239 ( .A(n10228), .B(n5684), .Z(n10241) );
  OR2 U6240 ( .A(n10242), .B(n10243), .Z(n10228) );
  OR2 U6241 ( .A(n10244), .B(n10245), .Z(n10243) );
  AN2 U6242 ( .A(n9968), .B(U156_Z_25), .Z(n10245) );
  AN2 U6243 ( .A(n10170), .B(U156_Z_20), .Z(n10244) );
  OR2 U6244 ( .A(n10038), .B(n10246), .Z(n10242) );
  AN2 U6245 ( .A(U61_DATA2_16), .B(n10147), .Z(n10246) );
  IV U6246 ( .A(n9223), .Z(n10239) );
  OR2 U6247 ( .A(n10247), .B(n10248), .Z(tx_data_out[53]) );
  AN2 U6248 ( .A(n9942), .B(n10249), .Z(n10248) );
  AN2 U6249 ( .A(n9929), .B(n9388), .Z(n10247) );
  OR2 U6250 ( .A(n10250), .B(n10251), .Z(n9388) );
  AN2 U6251 ( .A(n10252), .B(n10253), .Z(n10251) );
  AN2 U6252 ( .A(n10254), .B(U37_DATA1_51), .Z(n10250) );
  IV U6253 ( .A(n10252), .Z(n10254) );
  OR2 U6254 ( .A(n10255), .B(n10256), .Z(n10252) );
  AN2 U6255 ( .A(n9234), .B(n10257), .Z(n10256) );
  OR2 U6256 ( .A(n10258), .B(n9953), .Z(n10257) );
  AN2 U6257 ( .A(n10259), .B(n9955), .Z(n10258) );
  IV U6258 ( .A(n10249), .Z(n10259) );
  AN2 U6259 ( .A(n10260), .B(n10261), .Z(n10255) );
  OR2 U6260 ( .A(n10262), .B(n1934), .Z(n10261) );
  AN2 U6261 ( .A(n10249), .B(n5684), .Z(n10262) );
  OR2 U6262 ( .A(n10263), .B(n10264), .Z(n10249) );
  OR2 U6263 ( .A(n10265), .B(n10266), .Z(n10264) );
  AN2 U6264 ( .A(n9968), .B(U156_Z_24), .Z(n10266) );
  AN2 U6265 ( .A(n10170), .B(U156_Z_19), .Z(n10265) );
  OR2 U6266 ( .A(n10038), .B(n10267), .Z(n10263) );
  AN2 U6267 ( .A(U61_DATA2_15), .B(n10147), .Z(n10267) );
  IV U6268 ( .A(n9234), .Z(n10260) );
  OR2 U6269 ( .A(n10268), .B(n10269), .Z(tx_data_out[52]) );
  AN2 U6270 ( .A(n9942), .B(n10270), .Z(n10269) );
  AN2 U6271 ( .A(n9929), .B(n9399), .Z(n10268) );
  OR2 U6272 ( .A(n10271), .B(n10272), .Z(n9399) );
  AN2 U6273 ( .A(n10273), .B(n10274), .Z(n10272) );
  AN2 U6274 ( .A(n10275), .B(U37_DATA1_50), .Z(n10271) );
  IV U6275 ( .A(n10273), .Z(n10275) );
  OR2 U6276 ( .A(n10276), .B(n10277), .Z(n10273) );
  AN2 U6277 ( .A(n9333), .B(n10278), .Z(n10277) );
  OR2 U6278 ( .A(n10279), .B(n9953), .Z(n10278) );
  AN2 U6279 ( .A(n10280), .B(n9955), .Z(n10279) );
  IV U6280 ( .A(n10270), .Z(n10280) );
  AN2 U6281 ( .A(n10281), .B(n10282), .Z(n10276) );
  OR2 U6282 ( .A(n10283), .B(n1934), .Z(n10282) );
  AN2 U6283 ( .A(n10270), .B(n5684), .Z(n10283) );
  OR2 U6284 ( .A(n10284), .B(n10285), .Z(n10270) );
  OR2 U6285 ( .A(n10286), .B(n10215), .Z(n10285) );
  OR2 U6286 ( .A(n10287), .B(n10171), .Z(n10215) );
  AN2 U6287 ( .A(n10147), .B(n8775), .Z(n10171) );
  AN2 U6288 ( .A(n10288), .B(n10289), .Z(n8775) );
  AN2 U6289 ( .A(n5422), .B(n1712), .Z(n10289) );
  IV U6290 ( .A(n1654), .Z(n5422) );
  AN2 U6291 ( .A(n8777), .B(n10147), .Z(n10287) );
  AN2 U6292 ( .A(U154_Z_4), .B(n10290), .Z(n8777) );
  AN2 U6293 ( .A(n5420), .B(n1812), .Z(n10290) );
  IV U6294 ( .A(n1776), .Z(n5420) );
  AN2 U6295 ( .A(n10170), .B(n8669), .Z(n10286) );
  OR2 U6296 ( .A(n10195), .B(n10291), .Z(n10284) );
  AN2 U6297 ( .A(n9968), .B(n8668), .Z(n10291) );
  OR2 U6298 ( .A(n10292), .B(n4170), .Z(n8668) );
  AN2 U6299 ( .A(U162_DATA3_50), .B(n10092), .Z(n10292) );
  AN2 U6300 ( .A(n10293), .B(n10147), .Z(n10195) );
  OR2 U6301 ( .A(n10294), .B(n10124), .Z(n10147) );
  AN2 U6302 ( .A(n1927), .B(n10125), .Z(n10294) );
  OR2 U6303 ( .A(n8778), .B(n8774), .Z(n10293) );
  AN2 U6304 ( .A(n5421), .B(n10288), .Z(n8774) );
  IV U6305 ( .A(n1712), .Z(n5421) );
  AN2 U6306 ( .A(n5423), .B(n10223), .Z(n8778) );
  AN2 U6307 ( .A(n10288), .B(n10295), .Z(n10223) );
  AN2 U6308 ( .A(n1654), .B(n1712), .Z(n10295) );
  AN2 U6309 ( .A(U154_Z_4), .B(n10296), .Z(n10288) );
  AN2 U6310 ( .A(n1776), .B(n1812), .Z(n10296) );
  IV U6311 ( .A(n1603), .Z(n5423) );
  IV U6312 ( .A(n9333), .Z(n10281) );
  OR2 U6313 ( .A(n10297), .B(n10298), .Z(tx_data_out[51]) );
  AN2 U6314 ( .A(n9942), .B(n10299), .Z(n10298) );
  AN2 U6315 ( .A(n9929), .B(n9410), .Z(n10297) );
  OR2 U6316 ( .A(n10300), .B(n10301), .Z(n9410) );
  AN2 U6317 ( .A(n10302), .B(n10303), .Z(n10301) );
  AN2 U6318 ( .A(n10304), .B(U37_DATA1_49), .Z(n10300) );
  IV U6319 ( .A(n10302), .Z(n10304) );
  OR2 U6320 ( .A(n10305), .B(n10306), .Z(n10302) );
  AN2 U6321 ( .A(n9454), .B(n10307), .Z(n10306) );
  OR2 U6322 ( .A(n10308), .B(n9953), .Z(n10307) );
  AN2 U6323 ( .A(n10309), .B(n9955), .Z(n10308) );
  IV U6324 ( .A(n10299), .Z(n10309) );
  AN2 U6325 ( .A(n10310), .B(n10311), .Z(n10305) );
  OR2 U6326 ( .A(n10312), .B(n1934), .Z(n10311) );
  AN2 U6327 ( .A(n10299), .B(n5684), .Z(n10312) );
  OR2 U6328 ( .A(n10313), .B(n10314), .Z(n10299) );
  OR2 U6329 ( .A(n10315), .B(n10316), .Z(n10314) );
  AN2 U6330 ( .A(n10170), .B(U158_Z_9), .Z(n10316) );
  AN2 U6331 ( .A(n10317), .B(n10318), .Z(n10315) );
  OR2 U6332 ( .A(n8788), .B(n10319), .Z(n10317) );
  OR2 U6333 ( .A(n8785), .B(n10320), .Z(n10319) );
  AN2 U6334 ( .A(n9968), .B(U158_Z_11), .Z(n10313) );
  IV U6335 ( .A(n9454), .Z(n10310) );
  OR2 U6336 ( .A(n10321), .B(n10322), .Z(tx_data_out[50]) );
  AN2 U6337 ( .A(n9942), .B(n10323), .Z(n10322) );
  AN2 U6338 ( .A(n9929), .B(n9421), .Z(n10321) );
  OR2 U6339 ( .A(n10324), .B(n10325), .Z(n9421) );
  AN2 U6340 ( .A(n10326), .B(n10327), .Z(n10325) );
  AN2 U6341 ( .A(n10328), .B(U37_DATA1_48), .Z(n10324) );
  IV U6342 ( .A(n10326), .Z(n10328) );
  OR2 U6343 ( .A(n10329), .B(n10330), .Z(n10326) );
  AN2 U6344 ( .A(n9575), .B(n10331), .Z(n10330) );
  OR2 U6345 ( .A(n10332), .B(n9953), .Z(n10331) );
  AN2 U6346 ( .A(n10333), .B(n9955), .Z(n10332) );
  IV U6347 ( .A(n10323), .Z(n10333) );
  AN2 U6348 ( .A(n10334), .B(n10335), .Z(n10329) );
  OR2 U6349 ( .A(n10336), .B(n1934), .Z(n10335) );
  AN2 U6350 ( .A(n10323), .B(n5684), .Z(n10336) );
  OR2 U6351 ( .A(n10337), .B(n10338), .Z(n10323) );
  OR2 U6352 ( .A(n10339), .B(n10340), .Z(n10338) );
  AN2 U6353 ( .A(n9968), .B(U159_Z_7), .Z(n10340) );
  AN2 U6354 ( .A(n10170), .B(U159_Z_6), .Z(n10339) );
  AN2 U6355 ( .A(n10125), .B(n1906), .Z(n10170) );
  OR2 U6356 ( .A(n10341), .B(n10342), .Z(n10337) );
  AN2 U6357 ( .A(n10343), .B(n10318), .Z(n10342) );
  OR2 U6358 ( .A(n8789), .B(n10320), .Z(n10343) );
  AN2 U6359 ( .A(n10344), .B(n8792), .Z(n10320) );
  IV U6360 ( .A(n9575), .Z(n10334) );
  OR2 U6361 ( .A(n10345), .B(n10346), .Z(tx_data_out[5]) );
  OR2 U6362 ( .A(n10347), .B(n10348), .Z(n10346) );
  AN2 U6363 ( .A(n9928), .B(U157_Z_0), .Z(n10348) );
  AN2 U6364 ( .A(n9929), .B(n9999), .Z(n10347) );
  AN2 U6365 ( .A(n9930), .B(U40_DATA2_3), .Z(n10345) );
  OR2 U6366 ( .A(n10349), .B(n10350), .Z(tx_data_out[49]) );
  AN2 U6367 ( .A(n9942), .B(n10351), .Z(n10350) );
  AN2 U6368 ( .A(n9929), .B(n9432), .Z(n10349) );
  OR2 U6369 ( .A(n10352), .B(n10353), .Z(n9432) );
  AN2 U6370 ( .A(n10354), .B(n10355), .Z(n10353) );
  AN2 U6371 ( .A(n10356), .B(U37_DATA1_47), .Z(n10352) );
  IV U6372 ( .A(n10354), .Z(n10356) );
  OR2 U6373 ( .A(n10357), .B(n10358), .Z(n10354) );
  AN2 U6374 ( .A(n9696), .B(n10359), .Z(n10358) );
  OR2 U6375 ( .A(n10360), .B(n9953), .Z(n10359) );
  AN2 U6376 ( .A(n10361), .B(n9955), .Z(n10360) );
  IV U6377 ( .A(n10351), .Z(n10361) );
  AN2 U6378 ( .A(n10362), .B(n10363), .Z(n10357) );
  OR2 U6379 ( .A(n10364), .B(n1934), .Z(n10363) );
  AN2 U6380 ( .A(n10351), .B(n5684), .Z(n10364) );
  OR2 U6381 ( .A(n10365), .B(n10366), .Z(n10351) );
  OR2 U6382 ( .A(n10367), .B(n10368), .Z(n10366) );
  AN2 U6383 ( .A(n10369), .B(U157_Z_5), .Z(n10367) );
  OR2 U6384 ( .A(n10370), .B(n10371), .Z(n10365) );
  AN2 U6385 ( .A(n9968), .B(U156_Z_23), .Z(n10371) );
  IV U6386 ( .A(n9696), .Z(n10362) );
  OR2 U6387 ( .A(n10372), .B(n10373), .Z(tx_data_out[48]) );
  AN2 U6388 ( .A(n9942), .B(n10374), .Z(n10373) );
  AN2 U6389 ( .A(n9929), .B(n9443), .Z(n10372) );
  OR2 U6390 ( .A(n10375), .B(n10376), .Z(n9443) );
  AN2 U6391 ( .A(n10377), .B(n10378), .Z(n10376) );
  AN2 U6392 ( .A(n10379), .B(U37_DATA1_46), .Z(n10375) );
  IV U6393 ( .A(n10377), .Z(n10379) );
  OR2 U6394 ( .A(n10380), .B(n10381), .Z(n10377) );
  AN2 U6395 ( .A(n9817), .B(n10382), .Z(n10381) );
  OR2 U6396 ( .A(n10383), .B(n9953), .Z(n10382) );
  AN2 U6397 ( .A(n10384), .B(n9955), .Z(n10383) );
  IV U6398 ( .A(n10374), .Z(n10384) );
  AN2 U6399 ( .A(n10385), .B(n10386), .Z(n10380) );
  OR2 U6400 ( .A(n10387), .B(n1934), .Z(n10386) );
  AN2 U6401 ( .A(n10374), .B(n5684), .Z(n10387) );
  OR2 U6402 ( .A(n10388), .B(n10389), .Z(n10374) );
  OR2 U6403 ( .A(n10368), .B(n10390), .Z(n10389) );
  OR2 U6404 ( .A(n10391), .B(n10038), .Z(n10368) );
  AN2 U6405 ( .A(n10392), .B(n10318), .Z(n10391) );
  OR2 U6406 ( .A(n10393), .B(n10394), .Z(n10392) );
  AN2 U6407 ( .A(n8725), .B(n10395), .Z(n10394) );
  OR2 U6408 ( .A(n1337), .B(n5407), .Z(n10395) );
  IV U6409 ( .A(n1446), .Z(n5407) );
  AN2 U6410 ( .A(n10396), .B(n8792), .Z(n8725) );
  IV U6411 ( .A(n10344), .Z(n10396) );
  OR2 U6412 ( .A(n5406), .B(n5400), .Z(n10344) );
  IV U6413 ( .A(n1561), .Z(n5406) );
  AN2 U6414 ( .A(n10397), .B(n8792), .Z(n10393) );
  AN2 U6415 ( .A(n1617), .B(n10398), .Z(n8792) );
  AN2 U6416 ( .A(n1561), .B(n5400), .Z(n10397) );
  IV U6417 ( .A(n1498), .Z(n5400) );
  OR2 U6418 ( .A(n10399), .B(n10400), .Z(n10388) );
  AN2 U6419 ( .A(n10369), .B(U156_Z_18), .Z(n10400) );
  AN2 U6420 ( .A(n9968), .B(U156_Z_22), .Z(n10399) );
  IV U6421 ( .A(n9817), .Z(n10385) );
  AN2 U6422 ( .A(n10401), .B(n10402), .Z(n9817) );
  IV U6423 ( .A(n10403), .Z(n10402) );
  AN2 U6424 ( .A(n10404), .B(n10405), .Z(n10403) );
  OR2 U6425 ( .A(n10405), .B(n10404), .Z(n10401) );
  OR2 U6426 ( .A(n10406), .B(n10407), .Z(n10404) );
  AN2 U6427 ( .A(U37_DATA1_26), .B(n10408), .Z(n10407) );
  IV U6428 ( .A(U37_DATA1_7), .Z(n10408) );
  AN2 U6429 ( .A(U37_DATA1_7), .B(n10409), .Z(n10406) );
  OR2 U6430 ( .A(n10410), .B(n10411), .Z(n10405) );
  OR2 U6431 ( .A(n1934), .B(n10412), .Z(n10411) );
  AN2 U6432 ( .A(n10413), .B(U157_Z_2), .Z(n10412) );
  AN2 U6433 ( .A(U40_DATA2_7), .B(n10414), .Z(n10410) );
  OR2 U6434 ( .A(n10415), .B(n10416), .Z(tx_data_out[47]) );
  AN2 U6435 ( .A(n9942), .B(n10417), .Z(n10416) );
  AN2 U6436 ( .A(n9929), .B(n9465), .Z(n10415) );
  OR2 U6437 ( .A(n10418), .B(n10419), .Z(n9465) );
  AN2 U6438 ( .A(n10420), .B(n10421), .Z(n10419) );
  AN2 U6439 ( .A(n10422), .B(U37_DATA1_45), .Z(n10418) );
  IV U6440 ( .A(n10420), .Z(n10422) );
  OR2 U6441 ( .A(n10423), .B(n10424), .Z(n10420) );
  AN2 U6442 ( .A(n9835), .B(n10425), .Z(n10424) );
  OR2 U6443 ( .A(n10426), .B(n9953), .Z(n10425) );
  AN2 U6444 ( .A(n10427), .B(n9955), .Z(n10426) );
  IV U6445 ( .A(n10417), .Z(n10427) );
  AN2 U6446 ( .A(n10428), .B(n10429), .Z(n10423) );
  OR2 U6447 ( .A(n10430), .B(n1934), .Z(n10429) );
  AN2 U6448 ( .A(n10417), .B(n5684), .Z(n10430) );
  OR2 U6449 ( .A(n10431), .B(n10432), .Z(n10417) );
  OR2 U6450 ( .A(n10433), .B(n10434), .Z(n10432) );
  AN2 U6451 ( .A(n10369), .B(U156_Z_17), .Z(n10434) );
  AN2 U6452 ( .A(n9968), .B(U156_Z_21), .Z(n10433) );
  OR2 U6453 ( .A(n10038), .B(n10435), .Z(n10431) );
  AN2 U6454 ( .A(U61_DATA2_9), .B(n10318), .Z(n10435) );
  IV U6455 ( .A(n9835), .Z(n10428) );
  AN2 U6456 ( .A(n10436), .B(n10437), .Z(n9835) );
  IV U6457 ( .A(n10438), .Z(n10437) );
  AN2 U6458 ( .A(n10439), .B(n10440), .Z(n10438) );
  OR2 U6459 ( .A(n10440), .B(n10439), .Z(n10436) );
  OR2 U6460 ( .A(n10441), .B(n10442), .Z(n10439) );
  AN2 U6461 ( .A(U37_DATA1_25), .B(n10443), .Z(n10442) );
  IV U6462 ( .A(U37_DATA1_6), .Z(n10443) );
  AN2 U6463 ( .A(U37_DATA1_6), .B(n10444), .Z(n10441) );
  OR2 U6464 ( .A(n10445), .B(n10446), .Z(n10440) );
  OR2 U6465 ( .A(n1932), .B(n10447), .Z(n10446) );
  AN2 U6466 ( .A(n10413), .B(U156_Z_1), .Z(n10447) );
  AN2 U6467 ( .A(U40_DATA2_6), .B(n10414), .Z(n10445) );
  OR2 U6468 ( .A(n10448), .B(n10449), .Z(tx_data_out[46]) );
  AN2 U6469 ( .A(n9942), .B(n10450), .Z(n10449) );
  AN2 U6470 ( .A(n9929), .B(n9476), .Z(n10448) );
  OR2 U6471 ( .A(n10451), .B(n10452), .Z(n9476) );
  AN2 U6472 ( .A(n10453), .B(n10454), .Z(n10452) );
  AN2 U6473 ( .A(n10455), .B(U37_DATA1_44), .Z(n10451) );
  IV U6474 ( .A(n10453), .Z(n10455) );
  OR2 U6475 ( .A(n10456), .B(n10457), .Z(n10453) );
  AN2 U6476 ( .A(n9939), .B(n10458), .Z(n10457) );
  OR2 U6477 ( .A(n10459), .B(n9953), .Z(n10458) );
  AN2 U6478 ( .A(n10460), .B(n9955), .Z(n10459) );
  IV U6479 ( .A(n10450), .Z(n10460) );
  AN2 U6480 ( .A(n9948), .B(n10461), .Z(n10456) );
  OR2 U6481 ( .A(n10462), .B(n1934), .Z(n10461) );
  AN2 U6482 ( .A(n10450), .B(n5684), .Z(n10462) );
  OR2 U6483 ( .A(n10463), .B(n10464), .Z(n10450) );
  OR2 U6484 ( .A(n10465), .B(n10466), .Z(n10464) );
  AN2 U6485 ( .A(n10369), .B(U157_Z_4), .Z(n10466) );
  AN2 U6486 ( .A(n9968), .B(U156_Z_20), .Z(n10465) );
  OR2 U6487 ( .A(n10038), .B(n10467), .Z(n10463) );
  AN2 U6488 ( .A(U61_DATA2_8), .B(n10318), .Z(n10467) );
  IV U6489 ( .A(n9939), .Z(n9948) );
  AN2 U6490 ( .A(n10468), .B(n10469), .Z(n9939) );
  IV U6491 ( .A(n10470), .Z(n10469) );
  AN2 U6492 ( .A(n10471), .B(n10472), .Z(n10470) );
  OR2 U6493 ( .A(n10472), .B(n10471), .Z(n10468) );
  OR2 U6494 ( .A(n10473), .B(n10474), .Z(n10471) );
  AN2 U6495 ( .A(U37_DATA1_24), .B(n10475), .Z(n10474) );
  IV U6496 ( .A(U37_DATA1_5), .Z(n10475) );
  AN2 U6497 ( .A(U37_DATA1_5), .B(n10476), .Z(n10473) );
  OR2 U6498 ( .A(n10477), .B(n10478), .Z(n10472) );
  OR2 U6499 ( .A(n1934), .B(n10479), .Z(n10478) );
  AN2 U6500 ( .A(n10413), .B(U156_Z_0), .Z(n10479) );
  AN2 U6501 ( .A(U40_DATA2_5), .B(n10414), .Z(n10477) );
  OR2 U6502 ( .A(n10480), .B(n10481), .Z(tx_data_out[45]) );
  AN2 U6503 ( .A(n9942), .B(n10482), .Z(n10481) );
  AN2 U6504 ( .A(n9929), .B(n9487), .Z(n10480) );
  OR2 U6505 ( .A(n10483), .B(n10484), .Z(n9487) );
  AN2 U6506 ( .A(n10485), .B(n10486), .Z(n10484) );
  AN2 U6507 ( .A(n10487), .B(U37_DATA1_43), .Z(n10483) );
  IV U6508 ( .A(n10485), .Z(n10487) );
  OR2 U6509 ( .A(n10488), .B(n10489), .Z(n10485) );
  AN2 U6510 ( .A(n9974), .B(n10490), .Z(n10489) );
  OR2 U6511 ( .A(n10491), .B(n9953), .Z(n10490) );
  AN2 U6512 ( .A(n10492), .B(n9955), .Z(n10491) );
  IV U6513 ( .A(n10482), .Z(n10492) );
  AN2 U6514 ( .A(n9977), .B(n10493), .Z(n10488) );
  OR2 U6515 ( .A(n10494), .B(n1934), .Z(n10493) );
  AN2 U6516 ( .A(n10482), .B(n5684), .Z(n10494) );
  OR2 U6517 ( .A(n10495), .B(n10496), .Z(n10482) );
  OR2 U6518 ( .A(n10497), .B(n10390), .Z(n10496) );
  OR2 U6519 ( .A(n10498), .B(n10341), .Z(n10390) );
  AN2 U6520 ( .A(n10318), .B(n8786), .Z(n10341) );
  AN2 U6521 ( .A(n10499), .B(n10500), .Z(n8786) );
  AN2 U6522 ( .A(n5404), .B(n1728), .Z(n10500) );
  IV U6523 ( .A(n1666), .Z(n5404) );
  AN2 U6524 ( .A(n8788), .B(n10318), .Z(n10498) );
  AN2 U6525 ( .A(U154_Z_3), .B(n10501), .Z(n8788) );
  AN2 U6526 ( .A(n5402), .B(n1818), .Z(n10501) );
  IV U6527 ( .A(n1791), .Z(n5402) );
  AN2 U6528 ( .A(n10369), .B(U157_Z_3), .Z(n10497) );
  OR2 U6529 ( .A(n10370), .B(n10502), .Z(n10495) );
  AN2 U6530 ( .A(n9968), .B(U156_Z_19), .Z(n10502) );
  AN2 U6531 ( .A(n10503), .B(n10318), .Z(n10370) );
  OR2 U6532 ( .A(n10504), .B(n10124), .Z(n10318) );
  AN2 U6533 ( .A(n1924), .B(n10125), .Z(n10504) );
  OR2 U6534 ( .A(n8789), .B(n8785), .Z(n10503) );
  AN2 U6535 ( .A(n5403), .B(n10499), .Z(n8785) );
  IV U6536 ( .A(n1728), .Z(n5403) );
  AN2 U6537 ( .A(n5405), .B(n10398), .Z(n8789) );
  AN2 U6538 ( .A(n10499), .B(n10505), .Z(n10398) );
  AN2 U6539 ( .A(n1666), .B(n1728), .Z(n10505) );
  AN2 U6540 ( .A(U154_Z_3), .B(n10506), .Z(n10499) );
  AN2 U6541 ( .A(n1791), .B(n1818), .Z(n10506) );
  IV U6542 ( .A(n1617), .Z(n5405) );
  IV U6543 ( .A(n9974), .Z(n9977) );
  AN2 U6544 ( .A(n10507), .B(n10508), .Z(n9974) );
  IV U6545 ( .A(n10509), .Z(n10508) );
  AN2 U6546 ( .A(n10510), .B(n10511), .Z(n10509) );
  OR2 U6547 ( .A(n10511), .B(n10510), .Z(n10507) );
  OR2 U6548 ( .A(n10512), .B(n10513), .Z(n10510) );
  AN2 U6549 ( .A(U37_DATA1_23), .B(n10514), .Z(n10513) );
  IV U6550 ( .A(U37_DATA1_4), .Z(n10514) );
  AN2 U6551 ( .A(U37_DATA1_4), .B(n10515), .Z(n10512) );
  OR2 U6552 ( .A(n10516), .B(n10517), .Z(n10511) );
  OR2 U6553 ( .A(n1932), .B(n10518), .Z(n10517) );
  AN2 U6554 ( .A(n10413), .B(U157_Z_1), .Z(n10518) );
  AN2 U6555 ( .A(U40_DATA2_4), .B(n10414), .Z(n10516) );
  OR2 U6556 ( .A(n10519), .B(n10520), .Z(tx_data_out[44]) );
  AN2 U6557 ( .A(n9942), .B(n10521), .Z(n10520) );
  AN2 U6558 ( .A(n9929), .B(n9498), .Z(n10519) );
  OR2 U6559 ( .A(n10522), .B(n10523), .Z(n9498) );
  AN2 U6560 ( .A(n10524), .B(n10525), .Z(n10523) );
  AN2 U6561 ( .A(n10526), .B(U37_DATA1_42), .Z(n10522) );
  IV U6562 ( .A(n10524), .Z(n10526) );
  OR2 U6563 ( .A(n10527), .B(n10528), .Z(n10524) );
  AN2 U6564 ( .A(n9999), .B(n10529), .Z(n10528) );
  OR2 U6565 ( .A(n10530), .B(n9953), .Z(n10529) );
  AN2 U6566 ( .A(n10531), .B(n9955), .Z(n10530) );
  IV U6567 ( .A(n10521), .Z(n10531) );
  AN2 U6568 ( .A(n10002), .B(n10532), .Z(n10527) );
  OR2 U6569 ( .A(n10533), .B(n1934), .Z(n10532) );
  AN2 U6570 ( .A(n10521), .B(n5684), .Z(n10533) );
  OR2 U6571 ( .A(n10534), .B(n10535), .Z(n10521) );
  OR2 U6572 ( .A(n10536), .B(n10537), .Z(n10535) );
  AN2 U6573 ( .A(n9968), .B(n8669), .Z(n10537) );
  OR2 U6574 ( .A(n10538), .B(n4170), .Z(n8669) );
  AN2 U6575 ( .A(U162_DATA3_42), .B(n10092), .Z(n10538) );
  AN2 U6576 ( .A(n10539), .B(n10540), .Z(n10536) );
  OR2 U6577 ( .A(n8799), .B(n10541), .Z(n10539) );
  OR2 U6578 ( .A(n8796), .B(n10542), .Z(n10541) );
  AN2 U6579 ( .A(n10369), .B(U159_Z_5), .Z(n10534) );
  IV U6580 ( .A(n9999), .Z(n10002) );
  AN2 U6581 ( .A(n10543), .B(n10544), .Z(n9999) );
  IV U6582 ( .A(n10545), .Z(n10544) );
  AN2 U6583 ( .A(n10546), .B(n10547), .Z(n10545) );
  OR2 U6584 ( .A(n10547), .B(n10546), .Z(n10543) );
  OR2 U6585 ( .A(n10548), .B(n10549), .Z(n10546) );
  AN2 U6586 ( .A(U37_DATA1_22), .B(n10550), .Z(n10549) );
  IV U6587 ( .A(U37_DATA1_3), .Z(n10550) );
  AN2 U6588 ( .A(U37_DATA1_3), .B(n10551), .Z(n10548) );
  OR2 U6589 ( .A(n10552), .B(n10553), .Z(n10547) );
  OR2 U6590 ( .A(n1934), .B(n10554), .Z(n10553) );
  AN2 U6591 ( .A(n10413), .B(U157_Z_0), .Z(n10554) );
  AN2 U6592 ( .A(U40_DATA2_3), .B(n10414), .Z(n10552) );
  OR2 U6593 ( .A(n10555), .B(n10556), .Z(tx_data_out[43]) );
  AN2 U6594 ( .A(n9942), .B(n10557), .Z(n10556) );
  AN2 U6595 ( .A(n9929), .B(n9509), .Z(n10555) );
  OR2 U6596 ( .A(n10558), .B(n10559), .Z(n9509) );
  AN2 U6597 ( .A(n10560), .B(n10561), .Z(n10559) );
  AN2 U6598 ( .A(n10562), .B(U37_DATA1_41), .Z(n10558) );
  IV U6599 ( .A(n10560), .Z(n10562) );
  OR2 U6600 ( .A(n10563), .B(n10564), .Z(n10560) );
  AN2 U6601 ( .A(n10022), .B(n10565), .Z(n10564) );
  OR2 U6602 ( .A(n10566), .B(n9953), .Z(n10565) );
  AN2 U6603 ( .A(n10567), .B(n9955), .Z(n10566) );
  IV U6604 ( .A(n10557), .Z(n10567) );
  AN2 U6605 ( .A(n10025), .B(n10568), .Z(n10563) );
  OR2 U6606 ( .A(n10569), .B(n1934), .Z(n10568) );
  AN2 U6607 ( .A(n10557), .B(n5684), .Z(n10569) );
  OR2 U6608 ( .A(n10570), .B(n10571), .Z(n10557) );
  OR2 U6609 ( .A(n10572), .B(n10573), .Z(n10571) );
  AN2 U6610 ( .A(n10369), .B(U158_Z_8), .Z(n10573) );
  AN2 U6611 ( .A(n9968), .B(U158_Z_9), .Z(n10572) );
  OR2 U6612 ( .A(n10574), .B(n10575), .Z(n10570) );
  AN2 U6613 ( .A(n10576), .B(n10540), .Z(n10575) );
  OR2 U6614 ( .A(n8800), .B(n10542), .Z(n10576) );
  AN2 U6615 ( .A(n10577), .B(n8803), .Z(n10542) );
  IV U6616 ( .A(n10022), .Z(n10025) );
  OR2 U6617 ( .A(n10578), .B(n10579), .Z(tx_data_out[42]) );
  AN2 U6618 ( .A(n9942), .B(n10580), .Z(n10579) );
  AN2 U6619 ( .A(n9929), .B(n9520), .Z(n10578) );
  OR2 U6620 ( .A(n10581), .B(n10582), .Z(n9520) );
  AN2 U6621 ( .A(n10583), .B(n10584), .Z(n10582) );
  AN2 U6622 ( .A(n10585), .B(U37_DATA1_40), .Z(n10581) );
  IV U6623 ( .A(n10583), .Z(n10585) );
  OR2 U6624 ( .A(n10586), .B(n10587), .Z(n10583) );
  AN2 U6625 ( .A(n10053), .B(n10588), .Z(n10587) );
  OR2 U6626 ( .A(n10589), .B(n9953), .Z(n10588) );
  AN2 U6627 ( .A(n10590), .B(n9955), .Z(n10589) );
  IV U6628 ( .A(n10580), .Z(n10590) );
  AN2 U6629 ( .A(n10056), .B(n10591), .Z(n10586) );
  OR2 U6630 ( .A(n10592), .B(n1934), .Z(n10591) );
  AN2 U6631 ( .A(n10580), .B(n5684), .Z(n10592) );
  OR2 U6632 ( .A(n10593), .B(n10594), .Z(n10580) );
  OR2 U6633 ( .A(n10595), .B(n10596), .Z(n10594) );
  AN2 U6634 ( .A(n10369), .B(U159_Z_4), .Z(n10596) );
  AN2 U6635 ( .A(n10125), .B(n1900), .Z(n10369) );
  OR2 U6636 ( .A(n5247), .B(n8736), .Z(n1900) );
  OR2 U6637 ( .A(n5245), .B(n5246), .Z(n8736) );
  AN2 U6638 ( .A(n9968), .B(U159_Z_6), .Z(n10595) );
  OR2 U6639 ( .A(n10597), .B(n10598), .Z(n9968) );
  OR2 U6640 ( .A(n10599), .B(n8737), .Z(n10598) );
  OR2 U6641 ( .A(n99), .B(n5254), .Z(n10597) );
  OR2 U6642 ( .A(n10038), .B(n10600), .Z(n10593) );
  AN2 U6643 ( .A(n10601), .B(n10540), .Z(n10600) );
  OR2 U6644 ( .A(n10602), .B(n10603), .Z(n10601) );
  IV U6645 ( .A(n10053), .Z(n10056) );
  OR2 U6646 ( .A(n10604), .B(n10605), .Z(tx_data_out[41]) );
  AN2 U6647 ( .A(n9942), .B(n10606), .Z(n10605) );
  AN2 U6648 ( .A(n9929), .B(n9531), .Z(n10604) );
  OR2 U6649 ( .A(n10607), .B(n10608), .Z(n9531) );
  AN2 U6650 ( .A(n10609), .B(n10610), .Z(n10608) );
  AN2 U6651 ( .A(n10611), .B(U37_DATA1_39), .Z(n10607) );
  IV U6652 ( .A(n10609), .Z(n10611) );
  OR2 U6653 ( .A(n10612), .B(n10613), .Z(n10609) );
  AN2 U6654 ( .A(n10075), .B(n10614), .Z(n10613) );
  OR2 U6655 ( .A(n10615), .B(n9953), .Z(n10614) );
  AN2 U6656 ( .A(n10616), .B(n9955), .Z(n10615) );
  IV U6657 ( .A(n10606), .Z(n10616) );
  AN2 U6658 ( .A(n10078), .B(n10617), .Z(n10612) );
  OR2 U6659 ( .A(n10618), .B(n1934), .Z(n10617) );
  AN2 U6660 ( .A(n10606), .B(n5684), .Z(n10618) );
  OR2 U6661 ( .A(n10619), .B(n10620), .Z(n10606) );
  OR2 U6662 ( .A(n10621), .B(n10622), .Z(n10620) );
  OR2 U6663 ( .A(n10623), .B(n10624), .Z(n10619) );
  OR2 U6664 ( .A(n10625), .B(n10626), .Z(n10624) );
  AN2 U6665 ( .A(n10627), .B(U157_Z_5), .Z(n10626) );
  AN2 U6666 ( .A(n10603), .B(n10540), .Z(n10625) );
  OR2 U6667 ( .A(n10628), .B(n10629), .Z(n10603) );
  AN2 U6668 ( .A(n8727), .B(n10630), .Z(n10629) );
  OR2 U6669 ( .A(n1358), .B(n5388), .Z(n10630) );
  IV U6670 ( .A(n1456), .Z(n5388) );
  AN2 U6671 ( .A(n10631), .B(n8803), .Z(n8727) );
  IV U6672 ( .A(n10577), .Z(n10631) );
  OR2 U6673 ( .A(n5387), .B(n5380), .Z(n10577) );
  IV U6674 ( .A(n1568), .Z(n5387) );
  AN2 U6675 ( .A(n10632), .B(n8803), .Z(n10628) );
  AN2 U6676 ( .A(n1624), .B(n10633), .Z(n8803) );
  AN2 U6677 ( .A(n1568), .B(n5380), .Z(n10632) );
  IV U6678 ( .A(n1512), .Z(n5380) );
  AN2 U6679 ( .A(n10634), .B(U156_Z_16), .Z(n10623) );
  IV U6680 ( .A(n10075), .Z(n10078) );
  OR2 U6681 ( .A(n10635), .B(n10636), .Z(tx_data_out[40]) );
  AN2 U6682 ( .A(n9942), .B(n10637), .Z(n10636) );
  AN2 U6683 ( .A(n9929), .B(n9542), .Z(n10635) );
  OR2 U6684 ( .A(n10638), .B(n10639), .Z(n9542) );
  AN2 U6685 ( .A(n10640), .B(n10641), .Z(n10639) );
  AN2 U6686 ( .A(n10642), .B(U37_DATA1_38), .Z(n10638) );
  IV U6687 ( .A(n10640), .Z(n10642) );
  OR2 U6688 ( .A(n10643), .B(n10644), .Z(n10640) );
  AN2 U6689 ( .A(n10645), .B(n10104), .Z(n10644) );
  IV U6690 ( .A(U37_DATA1_57), .Z(n10104) );
  OR2 U6691 ( .A(n10646), .B(n1934), .Z(n10645) );
  AN2 U6692 ( .A(n10637), .B(n5684), .Z(n10646) );
  AN2 U6693 ( .A(U37_DATA1_57), .B(n10647), .Z(n10643) );
  OR2 U6694 ( .A(n10648), .B(n9953), .Z(n10647) );
  AN2 U6695 ( .A(n10649), .B(n9955), .Z(n10648) );
  IV U6696 ( .A(n10637), .Z(n10649) );
  OR2 U6697 ( .A(n10650), .B(n10651), .Z(n10637) );
  OR2 U6698 ( .A(n10652), .B(n10622), .Z(n10651) );
  AN2 U6699 ( .A(n10634), .B(U156_Z_15), .Z(n10652) );
  OR2 U6700 ( .A(n10653), .B(n10654), .Z(n10650) );
  AN2 U6701 ( .A(n10627), .B(U156_Z_18), .Z(n10654) );
  AN2 U6702 ( .A(U61_DATA2_2), .B(n10540), .Z(n10653) );
  OR2 U6703 ( .A(n10655), .B(n10656), .Z(tx_data_out[4]) );
  OR2 U6704 ( .A(n10657), .B(n10658), .Z(n10656) );
  AN2 U6705 ( .A(n9928), .B(U159_Z_1), .Z(n10658) );
  AN2 U6706 ( .A(n9929), .B(n10022), .Z(n10657) );
  AN2 U6707 ( .A(n10659), .B(n10660), .Z(n10022) );
  IV U6708 ( .A(n10661), .Z(n10660) );
  AN2 U6709 ( .A(n10662), .B(n10663), .Z(n10661) );
  OR2 U6710 ( .A(n10663), .B(n10662), .Z(n10659) );
  OR2 U6711 ( .A(n10664), .B(n10665), .Z(n10662) );
  AN2 U6712 ( .A(U37_DATA1_2), .B(n10666), .Z(n10665) );
  AN2 U6713 ( .A(U37_DATA1_21), .B(n10667), .Z(n10664) );
  IV U6714 ( .A(U37_DATA1_2), .Z(n10667) );
  OR2 U6715 ( .A(n10668), .B(n10669), .Z(n10663) );
  OR2 U6716 ( .A(n1932), .B(n10670), .Z(n10669) );
  AN2 U6717 ( .A(n10413), .B(U159_Z_1), .Z(n10670) );
  AN2 U6718 ( .A(U40_DATA2_2), .B(n10414), .Z(n10668) );
  AN2 U6719 ( .A(n9930), .B(U40_DATA2_2), .Z(n10655) );
  OR2 U6720 ( .A(n10671), .B(n10672), .Z(tx_data_out[39]) );
  AN2 U6721 ( .A(n9942), .B(n10673), .Z(n10672) );
  AN2 U6722 ( .A(n9929), .B(n9553), .Z(n10671) );
  OR2 U6723 ( .A(n10674), .B(n10675), .Z(n9553) );
  AN2 U6724 ( .A(n10676), .B(n10677), .Z(n10675) );
  AN2 U6725 ( .A(n10678), .B(U37_DATA1_37), .Z(n10674) );
  IV U6726 ( .A(n10676), .Z(n10678) );
  OR2 U6727 ( .A(n10679), .B(n10680), .Z(n10676) );
  AN2 U6728 ( .A(n10681), .B(n10139), .Z(n10680) );
  IV U6729 ( .A(U37_DATA1_56), .Z(n10139) );
  OR2 U6730 ( .A(n10682), .B(n1934), .Z(n10681) );
  AN2 U6731 ( .A(n10673), .B(n5684), .Z(n10682) );
  AN2 U6732 ( .A(U37_DATA1_56), .B(n10683), .Z(n10679) );
  OR2 U6733 ( .A(n10684), .B(n9953), .Z(n10683) );
  AN2 U6734 ( .A(n10685), .B(n9955), .Z(n10684) );
  IV U6735 ( .A(n10673), .Z(n10685) );
  OR2 U6736 ( .A(n10686), .B(n10687), .Z(n10673) );
  OR2 U6737 ( .A(n10688), .B(n10622), .Z(n10687) );
  OR2 U6738 ( .A(n10689), .B(n10038), .Z(n10622) );
  AN2 U6739 ( .A(n10634), .B(U156_Z_14), .Z(n10688) );
  OR2 U6740 ( .A(n10690), .B(n10691), .Z(n10686) );
  AN2 U6741 ( .A(n10627), .B(U156_Z_17), .Z(n10691) );
  AN2 U6742 ( .A(U61_DATA2_1), .B(n10540), .Z(n10690) );
  OR2 U6743 ( .A(n10692), .B(n10693), .Z(tx_data_out[38]) );
  AN2 U6744 ( .A(n9942), .B(n10694), .Z(n10693) );
  AN2 U6745 ( .A(n9929), .B(n9564), .Z(n10692) );
  OR2 U6746 ( .A(n10695), .B(n10696), .Z(n9564) );
  AN2 U6747 ( .A(n10697), .B(n10698), .Z(n10696) );
  AN2 U6748 ( .A(n10699), .B(U37_DATA1_36), .Z(n10695) );
  IV U6749 ( .A(n10697), .Z(n10699) );
  OR2 U6750 ( .A(n10700), .B(n10701), .Z(n10697) );
  AN2 U6751 ( .A(n10702), .B(n10156), .Z(n10701) );
  IV U6752 ( .A(U37_DATA1_55), .Z(n10156) );
  OR2 U6753 ( .A(n10703), .B(n1934), .Z(n10702) );
  AN2 U6754 ( .A(n10694), .B(n5684), .Z(n10703) );
  AN2 U6755 ( .A(U37_DATA1_55), .B(n10704), .Z(n10700) );
  OR2 U6756 ( .A(n10705), .B(n9953), .Z(n10704) );
  AN2 U6757 ( .A(n10706), .B(n9955), .Z(n10705) );
  IV U6758 ( .A(n10694), .Z(n10706) );
  OR2 U6759 ( .A(n10707), .B(n10708), .Z(n10694) );
  OR2 U6760 ( .A(n10709), .B(n10621), .Z(n10708) );
  OR2 U6761 ( .A(n10710), .B(n10574), .Z(n10621) );
  AN2 U6762 ( .A(n10540), .B(n8797), .Z(n10574) );
  AN2 U6763 ( .A(n10711), .B(n10712), .Z(n8797) );
  AN2 U6764 ( .A(n5385), .B(n1736), .Z(n10712) );
  IV U6765 ( .A(n1672), .Z(n5385) );
  AN2 U6766 ( .A(n8799), .B(n10540), .Z(n10710) );
  AN2 U6767 ( .A(U155_Z_1), .B(n10713), .Z(n8799) );
  AN2 U6768 ( .A(n5383), .B(n1821), .Z(n10713) );
  IV U6769 ( .A(n1798), .Z(n5383) );
  AN2 U6770 ( .A(n10634), .B(U156_Z_13), .Z(n10709) );
  OR2 U6771 ( .A(n10714), .B(n10715), .Z(n10707) );
  OR2 U6772 ( .A(n10689), .B(n10716), .Z(n10715) );
  AN2 U6773 ( .A(n10602), .B(n10540), .Z(n10716) );
  OR2 U6774 ( .A(n10717), .B(n10124), .Z(n10540) );
  AN2 U6775 ( .A(n2136), .B(n10718), .Z(n10124) );
  AN2 U6776 ( .A(n10125), .B(n8728), .Z(n10718) );
  AN2 U6777 ( .A(n1918), .B(n10125), .Z(n10717) );
  OR2 U6778 ( .A(n8800), .B(n8796), .Z(n10602) );
  AN2 U6779 ( .A(n5384), .B(n10711), .Z(n8796) );
  IV U6780 ( .A(n1736), .Z(n5384) );
  AN2 U6781 ( .A(n5386), .B(n10633), .Z(n8800) );
  AN2 U6782 ( .A(n10711), .B(n10719), .Z(n10633) );
  AN2 U6783 ( .A(n1672), .B(n1736), .Z(n10719) );
  AN2 U6784 ( .A(U155_Z_1), .B(n10720), .Z(n10711) );
  AN2 U6785 ( .A(n1798), .B(n1821), .Z(n10720) );
  IV U6786 ( .A(n1624), .Z(n5386) );
  AN2 U6787 ( .A(n10721), .B(n277), .Z(n10689) );
  AN2 U6788 ( .A(n10722), .B(n10125), .Z(n10721) );
  OR2 U6789 ( .A(n10599), .B(n1919), .Z(n10722) );
  AN2 U6790 ( .A(ALTERNATE_ENCODE), .B(n8728), .Z(n10599) );
  AN2 U6791 ( .A(n10627), .B(U157_Z_4), .Z(n10714) );
  OR2 U6792 ( .A(n10723), .B(n10724), .Z(tx_data_out[37]) );
  AN2 U6793 ( .A(n9942), .B(n10725), .Z(n10724) );
  AN2 U6794 ( .A(n9929), .B(n9586), .Z(n10723) );
  OR2 U6795 ( .A(n10726), .B(n10727), .Z(n9586) );
  AN2 U6796 ( .A(n10728), .B(n10729), .Z(n10727) );
  AN2 U6797 ( .A(n10730), .B(U37_DATA1_35), .Z(n10726) );
  IV U6798 ( .A(n10728), .Z(n10730) );
  OR2 U6799 ( .A(n10731), .B(n10732), .Z(n10728) );
  AN2 U6800 ( .A(n10733), .B(n10181), .Z(n10732) );
  IV U6801 ( .A(U37_DATA1_54), .Z(n10181) );
  OR2 U6802 ( .A(n10734), .B(n1934), .Z(n10733) );
  AN2 U6803 ( .A(n10725), .B(n5684), .Z(n10734) );
  AN2 U6804 ( .A(U37_DATA1_54), .B(n10735), .Z(n10731) );
  OR2 U6805 ( .A(n10736), .B(n9953), .Z(n10735) );
  AN2 U6806 ( .A(n10737), .B(n9955), .Z(n10736) );
  IV U6807 ( .A(n10725), .Z(n10737) );
  OR2 U6808 ( .A(n10738), .B(n10739), .Z(n10725) );
  OR2 U6809 ( .A(n10740), .B(n10741), .Z(n10739) );
  AN2 U6810 ( .A(n10634), .B(U156_Z_12), .Z(n10740) );
  OR2 U6811 ( .A(n10742), .B(n10743), .Z(n10738) );
  AN2 U6812 ( .A(n10627), .B(U157_Z_3), .Z(n10743) );
  AN2 U6813 ( .A(n10744), .B(n10745), .Z(n10742) );
  OR2 U6814 ( .A(n10746), .B(n10747), .Z(tx_data_out[36]) );
  AN2 U6815 ( .A(n9942), .B(n10748), .Z(n10747) );
  AN2 U6816 ( .A(n9929), .B(n9597), .Z(n10746) );
  OR2 U6817 ( .A(n10749), .B(n10750), .Z(n9597) );
  AN2 U6818 ( .A(n10751), .B(n10752), .Z(n10750) );
  AN2 U6819 ( .A(n10753), .B(U37_DATA1_34), .Z(n10749) );
  IV U6820 ( .A(n10751), .Z(n10753) );
  OR2 U6821 ( .A(n10754), .B(n10755), .Z(n10751) );
  AN2 U6822 ( .A(n10756), .B(n10203), .Z(n10755) );
  IV U6823 ( .A(U37_DATA1_53), .Z(n10203) );
  OR2 U6824 ( .A(n10757), .B(n1934), .Z(n10756) );
  AN2 U6825 ( .A(n10748), .B(n5684), .Z(n10757) );
  AN2 U6826 ( .A(U37_DATA1_53), .B(n10758), .Z(n10754) );
  OR2 U6827 ( .A(n10759), .B(n9953), .Z(n10758) );
  AN2 U6828 ( .A(n10760), .B(n9955), .Z(n10759) );
  IV U6829 ( .A(n10748), .Z(n10760) );
  OR2 U6830 ( .A(n10761), .B(n10762), .Z(n10748) );
  OR2 U6831 ( .A(n10763), .B(n10741), .Z(n10762) );
  OR2 U6832 ( .A(n10764), .B(n10765), .Z(n10741) );
  AN2 U6833 ( .A(n10766), .B(n273), .Z(n10765) );
  AN2 U6834 ( .A(n10767), .B(n10125), .Z(n10766) );
  AN2 U6835 ( .A(n10768), .B(n10744), .Z(n10764) );
  AN2 U6836 ( .A(n8814), .B(n10769), .Z(n10768) );
  IV U6837 ( .A(n10770), .Z(n10769) );
  AN2 U6838 ( .A(n10634), .B(n8670), .Z(n10763) );
  AN2 U6839 ( .A(n10125), .B(n10771), .Z(n10634) );
  OR2 U6840 ( .A(n10772), .B(n10773), .Z(n10761) );
  AN2 U6841 ( .A(n10627), .B(U159_Z_5), .Z(n10773) );
  OR2 U6842 ( .A(n8742), .B(n99), .Z(n10627) );
  AN2 U6843 ( .A(n10744), .B(n10774), .Z(n10772) );
  OR2 U6844 ( .A(n10775), .B(n10776), .Z(tx_data_out[35]) );
  OR2 U6845 ( .A(n10777), .B(n10778), .Z(n10776) );
  AN2 U6846 ( .A(n9930), .B(n10779), .Z(n10778) );
  AN2 U6847 ( .A(n9929), .B(n9608), .Z(n10777) );
  IV U6848 ( .A(n10780), .Z(n9608) );
  OR2 U6849 ( .A(n10781), .B(n10782), .Z(n10780) );
  AN2 U6850 ( .A(n10783), .B(n10784), .Z(n10782) );
  AN2 U6851 ( .A(n10785), .B(n10786), .Z(n10784) );
  OR2 U6852 ( .A(U37_DATA1_33), .B(n10232), .Z(n10786) );
  OR2 U6853 ( .A(U37_DATA1_52), .B(n10787), .Z(n10785) );
  IV U6854 ( .A(n10788), .Z(n10783) );
  AN2 U6855 ( .A(n10789), .B(n10788), .Z(n10781) );
  OR2 U6856 ( .A(n10790), .B(n10791), .Z(n10788) );
  OR2 U6857 ( .A(n1934), .B(n10792), .Z(n10791) );
  AN2 U6858 ( .A(n10414), .B(n10779), .Z(n10792) );
  OR2 U6859 ( .A(n10793), .B(n10794), .Z(n10779) );
  OR2 U6860 ( .A(n10795), .B(n10796), .Z(n10794) );
  AN2 U6861 ( .A(n8742), .B(U158_Z_8), .Z(n10795) );
  OR2 U6862 ( .A(n10797), .B(n10798), .Z(n10793) );
  AN2 U6863 ( .A(n10771), .B(U158_Z_6), .Z(n10798) );
  AN2 U6864 ( .A(n1914), .B(n10799), .Z(n10797) );
  OR2 U6865 ( .A(n8811), .B(n8808), .Z(n10799) );
  AN2 U6866 ( .A(n10413), .B(U158_Z_8), .Z(n10790) );
  OR2 U6867 ( .A(n10800), .B(n10801), .Z(n10789) );
  AN2 U6868 ( .A(U37_DATA1_33), .B(n10232), .Z(n10801) );
  IV U6869 ( .A(U37_DATA1_52), .Z(n10232) );
  AN2 U6870 ( .A(U37_DATA1_52), .B(n10787), .Z(n10800) );
  AN2 U6871 ( .A(n9928), .B(U158_Z_8), .Z(n10775) );
  OR2 U6872 ( .A(n10802), .B(n10803), .Z(tx_data_out[34]) );
  OR2 U6873 ( .A(n10804), .B(n10805), .Z(n10803) );
  AN2 U6874 ( .A(n9930), .B(n10806), .Z(n10805) );
  AN2 U6875 ( .A(n9929), .B(n9619), .Z(n10804) );
  IV U6876 ( .A(n10807), .Z(n9619) );
  OR2 U6877 ( .A(n10808), .B(n10809), .Z(n10807) );
  AN2 U6878 ( .A(n10810), .B(n10811), .Z(n10809) );
  AN2 U6879 ( .A(n10812), .B(n10813), .Z(n10811) );
  OR2 U6880 ( .A(U37_DATA1_32), .B(n10253), .Z(n10813) );
  OR2 U6881 ( .A(U37_DATA1_51), .B(n10814), .Z(n10812) );
  IV U6882 ( .A(n10815), .Z(n10810) );
  AN2 U6883 ( .A(n10816), .B(n10815), .Z(n10808) );
  OR2 U6884 ( .A(n10817), .B(n10818), .Z(n10815) );
  OR2 U6885 ( .A(n1934), .B(n10819), .Z(n10818) );
  AN2 U6886 ( .A(n10414), .B(n10806), .Z(n10819) );
  OR2 U6887 ( .A(n10820), .B(n10821), .Z(n10806) );
  OR2 U6888 ( .A(n10822), .B(n10796), .Z(n10821) );
  OR2 U6889 ( .A(n10823), .B(n10824), .Z(n10796) );
  OR2 U6890 ( .A(n8755), .B(n10825), .Z(n10824) );
  AN2 U6891 ( .A(n1914), .B(n10826), .Z(n10825) );
  OR2 U6892 ( .A(n10827), .B(n10828), .Z(n10826) );
  AN2 U6893 ( .A(n8815), .B(n10829), .Z(n10828) );
  OR2 U6894 ( .A(n1278), .B(n5368), .Z(n10829) );
  IV U6895 ( .A(n1371), .Z(n5368) );
  AN2 U6896 ( .A(n10770), .B(n8814), .Z(n8815) );
  AN2 U6897 ( .A(n1519), .B(n1462), .Z(n10770) );
  AN2 U6898 ( .A(n10830), .B(n8814), .Z(n10827) );
  AN2 U6899 ( .A(n1575), .B(n10831), .Z(n8814) );
  AN2 U6900 ( .A(n1519), .B(n5361), .Z(n10830) );
  IV U6901 ( .A(n1462), .Z(n5361) );
  AN2 U6902 ( .A(n273), .B(n10767), .Z(n10823) );
  AN2 U6903 ( .A(n8742), .B(U159_Z_4), .Z(n10822) );
  OR2 U6904 ( .A(n10832), .B(n10833), .Z(n10820) );
  AN2 U6905 ( .A(n10771), .B(U158_Z_5), .Z(n10833) );
  AN2 U6906 ( .A(n1914), .B(n10834), .Z(n10832) );
  OR2 U6907 ( .A(n8810), .B(n8807), .Z(n10834) );
  AN2 U6908 ( .A(n10413), .B(U159_Z_4), .Z(n10817) );
  OR2 U6909 ( .A(n10835), .B(n10836), .Z(n10816) );
  AN2 U6910 ( .A(U37_DATA1_32), .B(n10253), .Z(n10836) );
  IV U6911 ( .A(U37_DATA1_51), .Z(n10253) );
  AN2 U6912 ( .A(U37_DATA1_51), .B(n10814), .Z(n10835) );
  AN2 U6913 ( .A(n9928), .B(U159_Z_4), .Z(n10802) );
  OR2 U6914 ( .A(n10837), .B(n10838), .Z(tx_data_out[33]) );
  AN2 U6915 ( .A(n9942), .B(n10839), .Z(n10838) );
  AN2 U6916 ( .A(n9929), .B(n9630), .Z(n10837) );
  OR2 U6917 ( .A(n10840), .B(n10841), .Z(n9630) );
  AN2 U6918 ( .A(n10842), .B(n10843), .Z(n10841) );
  AN2 U6919 ( .A(n10844), .B(U37_DATA1_31), .Z(n10840) );
  IV U6920 ( .A(n10842), .Z(n10844) );
  OR2 U6921 ( .A(n10845), .B(n10846), .Z(n10842) );
  AN2 U6922 ( .A(n10847), .B(n10274), .Z(n10846) );
  IV U6923 ( .A(U37_DATA1_50), .Z(n10274) );
  OR2 U6924 ( .A(n10848), .B(n1934), .Z(n10847) );
  AN2 U6925 ( .A(n10839), .B(n5684), .Z(n10848) );
  AN2 U6926 ( .A(U37_DATA1_50), .B(n10849), .Z(n10845) );
  OR2 U6927 ( .A(n10850), .B(n9953), .Z(n10849) );
  AN2 U6928 ( .A(n10851), .B(n9955), .Z(n10850) );
  IV U6929 ( .A(n10839), .Z(n10851) );
  OR2 U6930 ( .A(n10852), .B(n10853), .Z(n10839) );
  OR2 U6931 ( .A(n10854), .B(n10855), .Z(n10853) );
  AN2 U6932 ( .A(n10856), .B(U156_Z_16), .Z(n10855) );
  AN2 U6933 ( .A(n10857), .B(U156_Z_11), .Z(n10854) );
  OR2 U6934 ( .A(n10038), .B(n10858), .Z(n10852) );
  AN2 U6935 ( .A(U52_DATA1_2), .B(n10744), .Z(n10858) );
  OR2 U6936 ( .A(n10859), .B(n10860), .Z(tx_data_out[32]) );
  AN2 U6937 ( .A(n9942), .B(n10861), .Z(n10860) );
  AN2 U6938 ( .A(n9929), .B(n9641), .Z(n10859) );
  OR2 U6939 ( .A(n10862), .B(n10863), .Z(n9641) );
  AN2 U6940 ( .A(n10864), .B(n10865), .Z(n10863) );
  AN2 U6941 ( .A(n10866), .B(U37_DATA1_30), .Z(n10862) );
  IV U6942 ( .A(n10864), .Z(n10866) );
  OR2 U6943 ( .A(n10867), .B(n10868), .Z(n10864) );
  AN2 U6944 ( .A(n10869), .B(n10303), .Z(n10868) );
  IV U6945 ( .A(U37_DATA1_49), .Z(n10303) );
  OR2 U6946 ( .A(n10870), .B(n1934), .Z(n10869) );
  AN2 U6947 ( .A(n10861), .B(n5684), .Z(n10870) );
  AN2 U6948 ( .A(U37_DATA1_49), .B(n10871), .Z(n10867) );
  OR2 U6949 ( .A(n10872), .B(n9953), .Z(n10871) );
  AN2 U6950 ( .A(n10873), .B(n9955), .Z(n10872) );
  IV U6951 ( .A(n10861), .Z(n10873) );
  OR2 U6952 ( .A(n10874), .B(n10875), .Z(n10861) );
  OR2 U6953 ( .A(n10876), .B(n10877), .Z(n10875) );
  AN2 U6954 ( .A(n10856), .B(U156_Z_15), .Z(n10877) );
  AN2 U6955 ( .A(n10857), .B(U156_Z_10), .Z(n10876) );
  OR2 U6956 ( .A(n10038), .B(n10878), .Z(n10874) );
  AN2 U6957 ( .A(U52_DATA1_1), .B(n10744), .Z(n10878) );
  OR2 U6958 ( .A(n10879), .B(n10880), .Z(tx_data_out[31]) );
  AN2 U6959 ( .A(n9942), .B(n10881), .Z(n10880) );
  AN2 U6960 ( .A(n9929), .B(n9652), .Z(n10879) );
  OR2 U6961 ( .A(n10882), .B(n10883), .Z(n9652) );
  AN2 U6962 ( .A(n10884), .B(n10885), .Z(n10883) );
  AN2 U6963 ( .A(n10886), .B(U37_DATA1_29), .Z(n10882) );
  IV U6964 ( .A(n10884), .Z(n10886) );
  OR2 U6965 ( .A(n10887), .B(n10888), .Z(n10884) );
  AN2 U6966 ( .A(n10889), .B(n10327), .Z(n10888) );
  IV U6967 ( .A(U37_DATA1_48), .Z(n10327) );
  OR2 U6968 ( .A(n10890), .B(n1934), .Z(n10889) );
  AN2 U6969 ( .A(n10881), .B(n5684), .Z(n10890) );
  AN2 U6970 ( .A(U37_DATA1_48), .B(n10891), .Z(n10887) );
  OR2 U6971 ( .A(n10892), .B(n9953), .Z(n10891) );
  AN2 U6972 ( .A(n10893), .B(n9955), .Z(n10892) );
  IV U6973 ( .A(n10881), .Z(n10893) );
  OR2 U6974 ( .A(n10894), .B(n10895), .Z(n10881) );
  OR2 U6975 ( .A(n10896), .B(n10897), .Z(n10895) );
  AN2 U6976 ( .A(n10857), .B(U156_Z_9), .Z(n10897) );
  AN2 U6977 ( .A(n10744), .B(n10898), .Z(n10896) );
  OR2 U6978 ( .A(n10774), .B(n10745), .Z(n10898) );
  OR2 U6979 ( .A(n8810), .B(n8808), .Z(n10745) );
  AN2 U6980 ( .A(n5364), .B(n10899), .Z(n8808) );
  IV U6981 ( .A(n1680), .Z(n5364) );
  AN2 U6982 ( .A(U154_Z_2), .B(n10900), .Z(n8810) );
  AN2 U6983 ( .A(n5363), .B(n1800), .Z(n10900) );
  IV U6984 ( .A(n1744), .Z(n5363) );
  OR2 U6985 ( .A(n8811), .B(n8807), .Z(n10774) );
  AN2 U6986 ( .A(n10899), .B(n10901), .Z(n8807) );
  AN2 U6987 ( .A(n5365), .B(n1680), .Z(n10901) );
  IV U6988 ( .A(n1630), .Z(n5365) );
  AN2 U6989 ( .A(n5366), .B(n10831), .Z(n8811) );
  AN2 U6990 ( .A(n10899), .B(n10902), .Z(n10831) );
  AN2 U6991 ( .A(n1630), .B(n1680), .Z(n10902) );
  AN2 U6992 ( .A(U154_Z_2), .B(n10903), .Z(n10899) );
  AN2 U6993 ( .A(n1744), .B(n1800), .Z(n10903) );
  IV U6994 ( .A(n1575), .Z(n5366) );
  AN2 U6995 ( .A(n10125), .B(n1914), .Z(n10744) );
  AN2 U6996 ( .A(n10856), .B(U156_Z_14), .Z(n10894) );
  OR2 U6997 ( .A(n10904), .B(n10905), .Z(tx_data_out[30]) );
  AN2 U6998 ( .A(n9942), .B(n10906), .Z(n10905) );
  AN2 U6999 ( .A(n9929), .B(n9663), .Z(n10904) );
  OR2 U7000 ( .A(n10907), .B(n10908), .Z(n9663) );
  AN2 U7001 ( .A(n10909), .B(n10910), .Z(n10908) );
  AN2 U7002 ( .A(n10911), .B(U37_DATA1_28), .Z(n10907) );
  IV U7003 ( .A(n10909), .Z(n10911) );
  OR2 U7004 ( .A(n10912), .B(n10913), .Z(n10909) );
  AN2 U7005 ( .A(n10914), .B(n10355), .Z(n10913) );
  IV U7006 ( .A(U37_DATA1_47), .Z(n10355) );
  OR2 U7007 ( .A(n10915), .B(n1934), .Z(n10914) );
  AN2 U7008 ( .A(n10906), .B(n5684), .Z(n10915) );
  AN2 U7009 ( .A(U37_DATA1_47), .B(n10916), .Z(n10912) );
  OR2 U7010 ( .A(n10917), .B(n9953), .Z(n10916) );
  AN2 U7011 ( .A(n10918), .B(n9955), .Z(n10917) );
  IV U7012 ( .A(n10906), .Z(n10918) );
  OR2 U7013 ( .A(n10919), .B(n10920), .Z(n10906) );
  OR2 U7014 ( .A(n10921), .B(n10922), .Z(n10920) );
  AN2 U7015 ( .A(n10857), .B(U156_Z_8), .Z(n10922) );
  AN2 U7016 ( .A(n10923), .B(n10924), .Z(n10921) );
  OR2 U7017 ( .A(n10925), .B(n10926), .Z(n10924) );
  AN2 U7018 ( .A(n10856), .B(U156_Z_13), .Z(n10919) );
  OR2 U7019 ( .A(n10927), .B(n10928), .Z(tx_data_out[3]) );
  OR2 U7020 ( .A(n10929), .B(n10930), .Z(n10928) );
  AN2 U7021 ( .A(n9928), .B(U158_Z_0), .Z(n10930) );
  AN2 U7022 ( .A(n9929), .B(n10053), .Z(n10929) );
  AN2 U7023 ( .A(n10931), .B(n10932), .Z(n10053) );
  IV U7024 ( .A(n10933), .Z(n10932) );
  AN2 U7025 ( .A(n10934), .B(n10935), .Z(n10933) );
  OR2 U7026 ( .A(n10935), .B(n10934), .Z(n10931) );
  OR2 U7027 ( .A(n10936), .B(n10937), .Z(n10934) );
  AN2 U7028 ( .A(U37_DATA1_1), .B(n10938), .Z(n10937) );
  AN2 U7029 ( .A(U37_DATA1_20), .B(n10939), .Z(n10936) );
  IV U7030 ( .A(U37_DATA1_1), .Z(n10939) );
  OR2 U7031 ( .A(n10940), .B(n10941), .Z(n10935) );
  OR2 U7032 ( .A(n1934), .B(n10942), .Z(n10941) );
  AN2 U7033 ( .A(n10413), .B(U158_Z_0), .Z(n10942) );
  AN2 U7034 ( .A(U40_DATA2_1), .B(n10414), .Z(n10940) );
  AN2 U7035 ( .A(n9930), .B(U40_DATA2_1), .Z(n10927) );
  OR2 U7036 ( .A(n10943), .B(n10944), .Z(tx_data_out[29]) );
  AN2 U7037 ( .A(n9942), .B(n10945), .Z(n10944) );
  AN2 U7038 ( .A(n9929), .B(n9674), .Z(n10943) );
  OR2 U7039 ( .A(n10946), .B(n10947), .Z(n9674) );
  AN2 U7040 ( .A(n10948), .B(n10949), .Z(n10947) );
  AN2 U7041 ( .A(n10950), .B(U37_DATA1_27), .Z(n10946) );
  IV U7042 ( .A(n10948), .Z(n10950) );
  OR2 U7043 ( .A(n10951), .B(n10952), .Z(n10948) );
  AN2 U7044 ( .A(n10953), .B(n10378), .Z(n10952) );
  IV U7045 ( .A(U37_DATA1_46), .Z(n10378) );
  OR2 U7046 ( .A(n10954), .B(n1934), .Z(n10953) );
  AN2 U7047 ( .A(n10945), .B(n5684), .Z(n10954) );
  AN2 U7048 ( .A(U37_DATA1_46), .B(n10955), .Z(n10951) );
  OR2 U7049 ( .A(n10956), .B(n9953), .Z(n10955) );
  AN2 U7050 ( .A(n10957), .B(n9955), .Z(n10956) );
  IV U7051 ( .A(n10945), .Z(n10957) );
  OR2 U7052 ( .A(n10958), .B(n10959), .Z(n10945) );
  OR2 U7053 ( .A(n10960), .B(n10961), .Z(n10959) );
  AN2 U7054 ( .A(n10857), .B(U156_Z_7), .Z(n10961) );
  AN2 U7055 ( .A(n10923), .B(n10962), .Z(n10960) );
  OR2 U7056 ( .A(n10925), .B(n10963), .Z(n10962) );
  AN2 U7057 ( .A(n10964), .B(n8826), .Z(n10925) );
  AN2 U7058 ( .A(n10856), .B(U156_Z_12), .Z(n10958) );
  OR2 U7059 ( .A(n10965), .B(n10966), .Z(tx_data_out[28]) );
  OR2 U7060 ( .A(n10967), .B(n10968), .Z(n10966) );
  AN2 U7061 ( .A(n9930), .B(n10969), .Z(n10968) );
  AN2 U7062 ( .A(n9929), .B(n9685), .Z(n10967) );
  IV U7063 ( .A(n10970), .Z(n9685) );
  OR2 U7064 ( .A(n10971), .B(n10972), .Z(n10970) );
  AN2 U7065 ( .A(n10973), .B(n10974), .Z(n10972) );
  AN2 U7066 ( .A(n10975), .B(n10976), .Z(n10974) );
  OR2 U7067 ( .A(U37_DATA1_26), .B(n10421), .Z(n10976) );
  OR2 U7068 ( .A(U37_DATA1_45), .B(n10409), .Z(n10975) );
  IV U7069 ( .A(n10977), .Z(n10973) );
  AN2 U7070 ( .A(n10978), .B(n10977), .Z(n10971) );
  OR2 U7071 ( .A(n10979), .B(n10980), .Z(n10977) );
  OR2 U7072 ( .A(n1934), .B(n10981), .Z(n10980) );
  AN2 U7073 ( .A(n10414), .B(n10969), .Z(n10981) );
  OR2 U7074 ( .A(n10982), .B(n10983), .Z(n10969) );
  OR2 U7075 ( .A(n10984), .B(n10985), .Z(n10983) );
  AN2 U7076 ( .A(n10986), .B(n8671), .Z(n10984) );
  OR2 U7077 ( .A(n10987), .B(n10988), .Z(n10982) );
  AN2 U7078 ( .A(n8735), .B(n8670), .Z(n10988) );
  AN2 U7079 ( .A(n10989), .B(n1898), .Z(n10987) );
  OR2 U7080 ( .A(n8823), .B(n8820), .Z(n10989) );
  AN2 U7081 ( .A(n10413), .B(n8670), .Z(n10979) );
  OR2 U7082 ( .A(n10990), .B(n10991), .Z(n10978) );
  AN2 U7083 ( .A(U37_DATA1_26), .B(n10421), .Z(n10991) );
  IV U7084 ( .A(U37_DATA1_45), .Z(n10421) );
  AN2 U7085 ( .A(U37_DATA1_45), .B(n10409), .Z(n10990) );
  IV U7086 ( .A(U37_DATA1_26), .Z(n10409) );
  AN2 U7087 ( .A(n9928), .B(n8670), .Z(n10965) );
  OR2 U7088 ( .A(n10992), .B(n4170), .Z(n8670) );
  AN2 U7089 ( .A(U162_DATA3_26), .B(n10092), .Z(n10992) );
  OR2 U7090 ( .A(n10993), .B(n10994), .Z(tx_data_out[27]) );
  OR2 U7091 ( .A(n10995), .B(n10996), .Z(n10994) );
  AN2 U7092 ( .A(n9930), .B(n10997), .Z(n10996) );
  AN2 U7093 ( .A(n9929), .B(n9707), .Z(n10995) );
  IV U7094 ( .A(n10998), .Z(n9707) );
  OR2 U7095 ( .A(n10999), .B(n11000), .Z(n10998) );
  AN2 U7096 ( .A(n11001), .B(n11002), .Z(n11000) );
  AN2 U7097 ( .A(n11003), .B(n11004), .Z(n11002) );
  OR2 U7098 ( .A(U37_DATA1_25), .B(n10454), .Z(n11004) );
  OR2 U7099 ( .A(U37_DATA1_44), .B(n10444), .Z(n11003) );
  IV U7100 ( .A(n11005), .Z(n11001) );
  AN2 U7101 ( .A(n11006), .B(n11005), .Z(n10999) );
  OR2 U7102 ( .A(n11007), .B(n11008), .Z(n11005) );
  OR2 U7103 ( .A(n1934), .B(n11009), .Z(n11008) );
  AN2 U7104 ( .A(n10414), .B(n10997), .Z(n11009) );
  OR2 U7105 ( .A(n11010), .B(n11011), .Z(n10997) );
  OR2 U7106 ( .A(n11012), .B(n10985), .Z(n11011) );
  OR2 U7107 ( .A(n11013), .B(n8755), .Z(n10985) );
  AN2 U7108 ( .A(n11014), .B(n1898), .Z(n11013) );
  OR2 U7109 ( .A(n11015), .B(n11016), .Z(n11014) );
  AN2 U7110 ( .A(n8827), .B(n11017), .Z(n11016) );
  OR2 U7111 ( .A(n1288), .B(n5350), .Z(n11017) );
  IV U7112 ( .A(n1384), .Z(n5350) );
  AN2 U7113 ( .A(n11018), .B(n8826), .Z(n8827) );
  IV U7114 ( .A(n10964), .Z(n11018) );
  OR2 U7115 ( .A(n5349), .B(n5343), .Z(n10964) );
  IV U7116 ( .A(n1526), .Z(n5349) );
  AN2 U7117 ( .A(n11019), .B(n8826), .Z(n11015) );
  AN2 U7118 ( .A(n1582), .B(n11020), .Z(n8826) );
  AN2 U7119 ( .A(n1526), .B(n5343), .Z(n11019) );
  IV U7120 ( .A(n1468), .Z(n5343) );
  AN2 U7121 ( .A(n8735), .B(U158_Z_6), .Z(n11012) );
  OR2 U7122 ( .A(n11021), .B(n11022), .Z(n11010) );
  AN2 U7123 ( .A(n10986), .B(U158_Z_3), .Z(n11022) );
  AN2 U7124 ( .A(n11023), .B(n1898), .Z(n11021) );
  OR2 U7125 ( .A(n8822), .B(n8819), .Z(n11023) );
  AN2 U7126 ( .A(n10413), .B(U158_Z_6), .Z(n11007) );
  OR2 U7127 ( .A(n11024), .B(n11025), .Z(n11006) );
  AN2 U7128 ( .A(U37_DATA1_25), .B(n10454), .Z(n11025) );
  IV U7129 ( .A(U37_DATA1_44), .Z(n10454) );
  AN2 U7130 ( .A(U37_DATA1_44), .B(n10444), .Z(n11024) );
  IV U7131 ( .A(U37_DATA1_25), .Z(n10444) );
  AN2 U7132 ( .A(n9928), .B(U158_Z_6), .Z(n10993) );
  OR2 U7133 ( .A(n11026), .B(n11027), .Z(tx_data_out[26]) );
  AN2 U7134 ( .A(n9942), .B(n11028), .Z(n11027) );
  AN2 U7135 ( .A(n9929), .B(n9718), .Z(n11026) );
  IV U7136 ( .A(n9956), .Z(n9718) );
  OR2 U7137 ( .A(n11029), .B(n11030), .Z(n9956) );
  AN2 U7138 ( .A(n11031), .B(n11032), .Z(n11030) );
  IV U7139 ( .A(n11033), .Z(n11029) );
  OR2 U7140 ( .A(n11032), .B(n11031), .Z(n11033) );
  OR2 U7141 ( .A(n11034), .B(n11035), .Z(n11031) );
  AN2 U7142 ( .A(U37_DATA1_24), .B(n10486), .Z(n11035) );
  IV U7143 ( .A(U37_DATA1_43), .Z(n10486) );
  AN2 U7144 ( .A(U37_DATA1_43), .B(n10476), .Z(n11034) );
  IV U7145 ( .A(U37_DATA1_24), .Z(n10476) );
  OR2 U7146 ( .A(n11036), .B(n1932), .Z(n11032) );
  AN2 U7147 ( .A(n11028), .B(n5684), .Z(n11036) );
  OR2 U7148 ( .A(n11037), .B(n11038), .Z(n11028) );
  OR2 U7149 ( .A(n11039), .B(n11040), .Z(n11038) );
  AN2 U7150 ( .A(n10856), .B(U158_Z_5), .Z(n11040) );
  AN2 U7151 ( .A(U54_DATA1_0), .B(n10923), .Z(n11039) );
  OR2 U7152 ( .A(n10038), .B(n11041), .Z(n11037) );
  AN2 U7153 ( .A(n10857), .B(U159_Z_3), .Z(n11041) );
  AN2 U7154 ( .A(n10125), .B(n10986), .Z(n10857) );
  OR2 U7155 ( .A(n11042), .B(n11043), .Z(tx_data_out[25]) );
  AN2 U7156 ( .A(n9942), .B(n11044), .Z(n11043) );
  AN2 U7157 ( .A(n9929), .B(n9729), .Z(n11042) );
  OR2 U7158 ( .A(n11045), .B(n11046), .Z(n9729) );
  AN2 U7159 ( .A(n11047), .B(n10515), .Z(n11046) );
  IV U7160 ( .A(U37_DATA1_23), .Z(n10515) );
  AN2 U7161 ( .A(n11048), .B(U37_DATA1_23), .Z(n11045) );
  IV U7162 ( .A(n11047), .Z(n11048) );
  OR2 U7163 ( .A(n11049), .B(n11050), .Z(n11047) );
  AN2 U7164 ( .A(n11051), .B(n10525), .Z(n11050) );
  IV U7165 ( .A(U37_DATA1_42), .Z(n10525) );
  OR2 U7166 ( .A(n11052), .B(n1934), .Z(n11051) );
  AN2 U7167 ( .A(n11044), .B(n5684), .Z(n11052) );
  AN2 U7168 ( .A(U37_DATA1_42), .B(n11053), .Z(n11049) );
  OR2 U7169 ( .A(n11054), .B(n9953), .Z(n11053) );
  AN2 U7170 ( .A(n11055), .B(n9955), .Z(n11054) );
  IV U7171 ( .A(n11044), .Z(n11055) );
  OR2 U7172 ( .A(n11056), .B(n11057), .Z(n11044) );
  OR2 U7173 ( .A(n11058), .B(n11059), .Z(n11057) );
  AN2 U7174 ( .A(n10856), .B(U156_Z_11), .Z(n11059) );
  AN2 U7175 ( .A(n11060), .B(U156_Z_6), .Z(n11058) );
  OR2 U7176 ( .A(n10038), .B(n11061), .Z(n11056) );
  AN2 U7177 ( .A(U55_DATA1_1), .B(n10923), .Z(n11061) );
  OR2 U7178 ( .A(n11062), .B(n11063), .Z(tx_data_out[24]) );
  AN2 U7179 ( .A(n9942), .B(n11064), .Z(n11063) );
  AN2 U7180 ( .A(n9929), .B(n9740), .Z(n11062) );
  OR2 U7181 ( .A(n11065), .B(n11066), .Z(n9740) );
  AN2 U7182 ( .A(n11067), .B(n10551), .Z(n11066) );
  IV U7183 ( .A(U37_DATA1_22), .Z(n10551) );
  AN2 U7184 ( .A(n11068), .B(U37_DATA1_22), .Z(n11065) );
  IV U7185 ( .A(n11067), .Z(n11068) );
  OR2 U7186 ( .A(n11069), .B(n11070), .Z(n11067) );
  AN2 U7187 ( .A(n11071), .B(n10561), .Z(n11070) );
  IV U7188 ( .A(U37_DATA1_41), .Z(n10561) );
  OR2 U7189 ( .A(n11072), .B(n1934), .Z(n11071) );
  AN2 U7190 ( .A(n11064), .B(n5684), .Z(n11072) );
  AN2 U7191 ( .A(U37_DATA1_41), .B(n11073), .Z(n11069) );
  OR2 U7192 ( .A(n11074), .B(n9953), .Z(n11073) );
  AN2 U7193 ( .A(n11075), .B(n9955), .Z(n11074) );
  IV U7194 ( .A(n11064), .Z(n11075) );
  OR2 U7195 ( .A(n11076), .B(n11077), .Z(n11064) );
  OR2 U7196 ( .A(n11078), .B(n11079), .Z(n11077) );
  AN2 U7197 ( .A(n11060), .B(U156_Z_5), .Z(n11079) );
  AN2 U7198 ( .A(n10923), .B(n11080), .Z(n11078) );
  OR2 U7199 ( .A(n10926), .B(n10963), .Z(n11080) );
  OR2 U7200 ( .A(n8823), .B(n8819), .Z(n10963) );
  AN2 U7201 ( .A(n11081), .B(n11082), .Z(n8819) );
  AN2 U7202 ( .A(n5347), .B(n1688), .Z(n11082) );
  IV U7203 ( .A(n1636), .Z(n5347) );
  AN2 U7204 ( .A(n5348), .B(n11020), .Z(n8823) );
  AN2 U7205 ( .A(n11081), .B(n11083), .Z(n11020) );
  AN2 U7206 ( .A(n1636), .B(n1688), .Z(n11083) );
  IV U7207 ( .A(n1582), .Z(n5348) );
  OR2 U7208 ( .A(n8822), .B(n8820), .Z(n10926) );
  AN2 U7209 ( .A(n5346), .B(n11081), .Z(n8820) );
  AN2 U7210 ( .A(U154_Z_1), .B(n11084), .Z(n11081) );
  AN2 U7211 ( .A(n1752), .B(n1803), .Z(n11084) );
  IV U7212 ( .A(n1688), .Z(n5346) );
  AN2 U7213 ( .A(U154_Z_1), .B(n11085), .Z(n8822) );
  AN2 U7214 ( .A(n5345), .B(n1803), .Z(n11085) );
  IV U7215 ( .A(n1752), .Z(n5345) );
  AN2 U7216 ( .A(n10125), .B(n1898), .Z(n10923) );
  OR2 U7217 ( .A(n8734), .B(n11086), .Z(n1898) );
  AN2 U7218 ( .A(n10856), .B(U156_Z_10), .Z(n11076) );
  OR2 U7219 ( .A(n11087), .B(n11088), .Z(tx_data_out[23]) );
  AN2 U7220 ( .A(n9942), .B(n11089), .Z(n11088) );
  AN2 U7221 ( .A(n9929), .B(n9751), .Z(n11087) );
  OR2 U7222 ( .A(n11090), .B(n11091), .Z(n9751) );
  AN2 U7223 ( .A(n11092), .B(n10666), .Z(n11091) );
  IV U7224 ( .A(U37_DATA1_21), .Z(n10666) );
  AN2 U7225 ( .A(n11093), .B(U37_DATA1_21), .Z(n11090) );
  IV U7226 ( .A(n11092), .Z(n11093) );
  OR2 U7227 ( .A(n11094), .B(n11095), .Z(n11092) );
  AN2 U7228 ( .A(n11096), .B(n10584), .Z(n11095) );
  IV U7229 ( .A(U37_DATA1_40), .Z(n10584) );
  OR2 U7230 ( .A(n11097), .B(n1934), .Z(n11096) );
  AN2 U7231 ( .A(n11089), .B(n5684), .Z(n11097) );
  AN2 U7232 ( .A(U37_DATA1_40), .B(n11098), .Z(n11094) );
  OR2 U7233 ( .A(n11099), .B(n9953), .Z(n11098) );
  AN2 U7234 ( .A(n11100), .B(n9955), .Z(n11099) );
  IV U7235 ( .A(n11089), .Z(n11100) );
  OR2 U7236 ( .A(n11101), .B(n11102), .Z(n11089) );
  OR2 U7237 ( .A(n11103), .B(n11104), .Z(n11102) );
  AN2 U7238 ( .A(n11060), .B(U156_Z_4), .Z(n11104) );
  AN2 U7239 ( .A(n11105), .B(n11106), .Z(n11103) );
  OR2 U7240 ( .A(n11107), .B(n11108), .Z(n11106) );
  AN2 U7241 ( .A(n10856), .B(U156_Z_9), .Z(n11101) );
  OR2 U7242 ( .A(n11109), .B(n11110), .Z(tx_data_out[22]) );
  AN2 U7243 ( .A(n9942), .B(n11111), .Z(n11110) );
  AN2 U7244 ( .A(n9929), .B(n9762), .Z(n11109) );
  OR2 U7245 ( .A(n11112), .B(n11113), .Z(n9762) );
  AN2 U7246 ( .A(n11114), .B(n10938), .Z(n11113) );
  IV U7247 ( .A(U37_DATA1_20), .Z(n10938) );
  AN2 U7248 ( .A(n11115), .B(U37_DATA1_20), .Z(n11112) );
  IV U7249 ( .A(n11114), .Z(n11115) );
  OR2 U7250 ( .A(n11116), .B(n11117), .Z(n11114) );
  AN2 U7251 ( .A(n11118), .B(n10610), .Z(n11117) );
  IV U7252 ( .A(U37_DATA1_39), .Z(n10610) );
  OR2 U7253 ( .A(n11119), .B(n1934), .Z(n11118) );
  AN2 U7254 ( .A(n11111), .B(n5684), .Z(n11119) );
  AN2 U7255 ( .A(U37_DATA1_39), .B(n11120), .Z(n11116) );
  OR2 U7256 ( .A(n11121), .B(n9953), .Z(n11120) );
  AN2 U7257 ( .A(n11122), .B(n9955), .Z(n11121) );
  IV U7258 ( .A(n11111), .Z(n11122) );
  OR2 U7259 ( .A(n11123), .B(n11124), .Z(n11111) );
  OR2 U7260 ( .A(n11125), .B(n11126), .Z(n11124) );
  AN2 U7261 ( .A(n11060), .B(U156_Z_3), .Z(n11126) );
  AN2 U7262 ( .A(n11105), .B(n11127), .Z(n11125) );
  OR2 U7263 ( .A(n11107), .B(n11128), .Z(n11127) );
  AN2 U7264 ( .A(n11129), .B(n8838), .Z(n11107) );
  AN2 U7265 ( .A(n10856), .B(U156_Z_8), .Z(n11123) );
  OR2 U7266 ( .A(n11130), .B(n11131), .Z(tx_data_out[21]) );
  OR2 U7267 ( .A(n11132), .B(n11133), .Z(n11131) );
  AN2 U7268 ( .A(n9930), .B(n11134), .Z(n11133) );
  AN2 U7269 ( .A(n9929), .B(n9773), .Z(n11132) );
  IV U7270 ( .A(n10084), .Z(n9773) );
  OR2 U7271 ( .A(n11135), .B(n11136), .Z(n10084) );
  AN2 U7272 ( .A(n11137), .B(n11138), .Z(n11136) );
  IV U7273 ( .A(n11139), .Z(n11135) );
  OR2 U7274 ( .A(n11138), .B(n11137), .Z(n11139) );
  OR2 U7275 ( .A(n11140), .B(n11141), .Z(n11137) );
  AN2 U7276 ( .A(U37_DATA1_19), .B(n10641), .Z(n11141) );
  IV U7277 ( .A(U37_DATA1_38), .Z(n10641) );
  AN2 U7278 ( .A(U37_DATA1_38), .B(n11142), .Z(n11140) );
  OR2 U7279 ( .A(n11143), .B(n11144), .Z(n11138) );
  OR2 U7280 ( .A(n1934), .B(n11145), .Z(n11144) );
  AN2 U7281 ( .A(n10414), .B(n11134), .Z(n11145) );
  OR2 U7282 ( .A(n11146), .B(n11147), .Z(n11134) );
  OR2 U7283 ( .A(n11148), .B(n11149), .Z(n11147) );
  AN2 U7284 ( .A(n1910), .B(U156_Z_2), .Z(n11148) );
  OR2 U7285 ( .A(n11150), .B(n11151), .Z(n11146) );
  AN2 U7286 ( .A(n8735), .B(U156_Z_7), .Z(n11151) );
  AN2 U7287 ( .A(n11152), .B(n11086), .Z(n11150) );
  OR2 U7288 ( .A(n8835), .B(n8832), .Z(n11152) );
  AN2 U7289 ( .A(n10413), .B(U156_Z_7), .Z(n11143) );
  AN2 U7290 ( .A(n9928), .B(U156_Z_7), .Z(n11130) );
  OR2 U7291 ( .A(n11153), .B(n11154), .Z(tx_data_out[20]) );
  OR2 U7292 ( .A(n11155), .B(n11156), .Z(n11154) );
  AN2 U7293 ( .A(n9930), .B(n11157), .Z(n11156) );
  AN2 U7294 ( .A(n9929), .B(n9784), .Z(n11155) );
  AN2 U7295 ( .A(n11158), .B(n11159), .Z(n9784) );
  IV U7296 ( .A(n11160), .Z(n11159) );
  AN2 U7297 ( .A(n11161), .B(n11162), .Z(n11160) );
  OR2 U7298 ( .A(n11162), .B(n11161), .Z(n11158) );
  OR2 U7299 ( .A(n11163), .B(n11164), .Z(n11161) );
  AN2 U7300 ( .A(U37_DATA1_18), .B(n10677), .Z(n11164) );
  IV U7301 ( .A(U37_DATA1_37), .Z(n10677) );
  AN2 U7302 ( .A(U37_DATA1_37), .B(n11165), .Z(n11163) );
  IV U7303 ( .A(U37_DATA1_18), .Z(n11165) );
  OR2 U7304 ( .A(n11166), .B(n11167), .Z(n11162) );
  OR2 U7305 ( .A(n1934), .B(n11168), .Z(n11167) );
  AN2 U7306 ( .A(n10414), .B(n11157), .Z(n11168) );
  OR2 U7307 ( .A(n11169), .B(n11170), .Z(n11157) );
  OR2 U7308 ( .A(n11171), .B(n11149), .Z(n11170) );
  OR2 U7309 ( .A(n11172), .B(n8755), .Z(n11149) );
  AN2 U7310 ( .A(n11173), .B(n11086), .Z(n11172) );
  OR2 U7311 ( .A(n11174), .B(n11175), .Z(n11173) );
  AN2 U7312 ( .A(n8839), .B(n11176), .Z(n11175) );
  OR2 U7313 ( .A(n1308), .B(n5332), .Z(n11176) );
  IV U7314 ( .A(n1410), .Z(n5332) );
  AN2 U7315 ( .A(n11177), .B(n8838), .Z(n8839) );
  IV U7316 ( .A(n11129), .Z(n11177) );
  OR2 U7317 ( .A(n5331), .B(n5325), .Z(n11129) );
  IV U7318 ( .A(n1540), .Z(n5331) );
  AN2 U7319 ( .A(n11178), .B(n8838), .Z(n11174) );
  AN2 U7320 ( .A(n1596), .B(n11179), .Z(n8838) );
  AN2 U7321 ( .A(n1540), .B(n5325), .Z(n11178) );
  IV U7322 ( .A(n1480), .Z(n5325) );
  AN2 U7323 ( .A(n1910), .B(n8672), .Z(n11171) );
  OR2 U7324 ( .A(n11180), .B(n11181), .Z(n11169) );
  AN2 U7325 ( .A(n8735), .B(n8671), .Z(n11181) );
  AN2 U7326 ( .A(n11182), .B(n11086), .Z(n11180) );
  OR2 U7327 ( .A(n8834), .B(n8831), .Z(n11182) );
  AN2 U7328 ( .A(n10413), .B(n8671), .Z(n11166) );
  AN2 U7329 ( .A(n9928), .B(n8671), .Z(n11153) );
  OR2 U7330 ( .A(n11183), .B(n4170), .Z(n8671) );
  AN2 U7331 ( .A(U162_DATA3_18), .B(n10092), .Z(n11183) );
  OR2 U7332 ( .A(n11184), .B(n11185), .Z(tx_data_out[2]) );
  AN2 U7333 ( .A(n9942), .B(n11186), .Z(n11185) );
  AN2 U7334 ( .A(n9929), .B(n10075), .Z(n11184) );
  AN2 U7335 ( .A(n11187), .B(n11188), .Z(n10075) );
  IV U7336 ( .A(n11189), .Z(n11188) );
  AN2 U7337 ( .A(n11190), .B(n11191), .Z(n11189) );
  OR2 U7338 ( .A(n11191), .B(n11190), .Z(n11187) );
  OR2 U7339 ( .A(n11192), .B(n11193), .Z(n11190) );
  AN2 U7340 ( .A(U37_DATA1_0), .B(n11142), .Z(n11193) );
  IV U7341 ( .A(U37_DATA1_19), .Z(n11142) );
  AN2 U7342 ( .A(U37_DATA1_19), .B(n11194), .Z(n11192) );
  IV U7343 ( .A(U37_DATA1_0), .Z(n11194) );
  OR2 U7344 ( .A(n11195), .B(n1932), .Z(n11191) );
  AN2 U7345 ( .A(n11186), .B(n5684), .Z(n11195) );
  OR2 U7346 ( .A(n11196), .B(n11197), .Z(n11186) );
  AN2 U7347 ( .A(n99), .B(U159_Z_0), .Z(n11197) );
  AN2 U7348 ( .A(U40_DATA2_0), .B(n10125), .Z(n11196) );
  OR2 U7349 ( .A(n11198), .B(n11199), .Z(tx_data_out[19]) );
  AN2 U7350 ( .A(n9942), .B(n11200), .Z(n11199) );
  AN2 U7351 ( .A(n9929), .B(n9795), .Z(n11198) );
  OR2 U7352 ( .A(n11201), .B(n11202), .Z(n9795) );
  AN2 U7353 ( .A(n11203), .B(n11204), .Z(n11202) );
  IV U7354 ( .A(U37_DATA1_17), .Z(n11204) );
  AN2 U7355 ( .A(n11205), .B(U37_DATA1_17), .Z(n11201) );
  IV U7356 ( .A(n11203), .Z(n11205) );
  OR2 U7357 ( .A(n11206), .B(n11207), .Z(n11203) );
  AN2 U7358 ( .A(n11208), .B(n10698), .Z(n11207) );
  IV U7359 ( .A(U37_DATA1_36), .Z(n10698) );
  OR2 U7360 ( .A(n11209), .B(n1934), .Z(n11208) );
  AN2 U7361 ( .A(n11200), .B(n5684), .Z(n11209) );
  AN2 U7362 ( .A(U37_DATA1_36), .B(n11210), .Z(n11206) );
  OR2 U7363 ( .A(n11211), .B(n9953), .Z(n11210) );
  AN2 U7364 ( .A(n11212), .B(n9955), .Z(n11211) );
  IV U7365 ( .A(n11200), .Z(n11212) );
  OR2 U7366 ( .A(n11213), .B(n11214), .Z(n11200) );
  OR2 U7367 ( .A(n11215), .B(n11216), .Z(n11214) );
  AN2 U7368 ( .A(n10856), .B(U158_Z_3), .Z(n11216) );
  AN2 U7369 ( .A(U57_DATA1_1), .B(n11105), .Z(n11215) );
  OR2 U7370 ( .A(n10038), .B(n11217), .Z(n11213) );
  AN2 U7371 ( .A(n11060), .B(U158_Z_1), .Z(n11217) );
  OR2 U7372 ( .A(n11218), .B(n11219), .Z(tx_data_out[18]) );
  AN2 U7373 ( .A(n9942), .B(n11220), .Z(n11219) );
  AN2 U7374 ( .A(n9929), .B(n9806), .Z(n11218) );
  OR2 U7375 ( .A(n11221), .B(n11222), .Z(n9806) );
  AN2 U7376 ( .A(n11223), .B(n11224), .Z(n11222) );
  IV U7377 ( .A(U37_DATA1_16), .Z(n11224) );
  AN2 U7378 ( .A(n11225), .B(U37_DATA1_16), .Z(n11221) );
  IV U7379 ( .A(n11223), .Z(n11225) );
  OR2 U7380 ( .A(n11226), .B(n11227), .Z(n11223) );
  AN2 U7381 ( .A(n11228), .B(n10729), .Z(n11227) );
  IV U7382 ( .A(U37_DATA1_35), .Z(n10729) );
  OR2 U7383 ( .A(n11229), .B(n1934), .Z(n11228) );
  AN2 U7384 ( .A(n11220), .B(n5684), .Z(n11229) );
  AN2 U7385 ( .A(U37_DATA1_35), .B(n11230), .Z(n11226) );
  OR2 U7386 ( .A(n11231), .B(n9953), .Z(n11230) );
  AN2 U7387 ( .A(n11232), .B(n9955), .Z(n11231) );
  IV U7388 ( .A(n11220), .Z(n11232) );
  OR2 U7389 ( .A(n11233), .B(n11234), .Z(n11220) );
  OR2 U7390 ( .A(n11235), .B(n11236), .Z(n11234) );
  AN2 U7391 ( .A(n10856), .B(U159_Z_3), .Z(n11236) );
  AN2 U7392 ( .A(U57_DATA1_0), .B(n11105), .Z(n11235) );
  OR2 U7393 ( .A(n10038), .B(n11237), .Z(n11233) );
  AN2 U7394 ( .A(n11060), .B(U159_Z_2), .Z(n11237) );
  AN2 U7395 ( .A(n10125), .B(n1910), .Z(n11060) );
  OR2 U7396 ( .A(n11238), .B(n11239), .Z(tx_data_out[17]) );
  AN2 U7397 ( .A(n9942), .B(n11240), .Z(n11239) );
  AN2 U7398 ( .A(n9929), .B(n9200), .Z(n11238) );
  OR2 U7399 ( .A(n11241), .B(n11242), .Z(n9200) );
  AN2 U7400 ( .A(n11243), .B(n11244), .Z(n11242) );
  IV U7401 ( .A(U37_DATA1_15), .Z(n11244) );
  AN2 U7402 ( .A(n11245), .B(U37_DATA1_15), .Z(n11241) );
  IV U7403 ( .A(n11243), .Z(n11245) );
  OR2 U7404 ( .A(n11246), .B(n11247), .Z(n11243) );
  AN2 U7405 ( .A(n11248), .B(n10752), .Z(n11247) );
  IV U7406 ( .A(U37_DATA1_34), .Z(n10752) );
  OR2 U7407 ( .A(n11249), .B(n1934), .Z(n11248) );
  AN2 U7408 ( .A(n11240), .B(n5684), .Z(n11249) );
  AN2 U7409 ( .A(U37_DATA1_34), .B(n11250), .Z(n11246) );
  OR2 U7410 ( .A(n11251), .B(n9953), .Z(n11250) );
  AN2 U7411 ( .A(n11252), .B(n9955), .Z(n11251) );
  IV U7412 ( .A(n11240), .Z(n11252) );
  OR2 U7413 ( .A(n11253), .B(n11254), .Z(n11240) );
  OR2 U7414 ( .A(n11255), .B(n11256), .Z(n11254) );
  AN2 U7415 ( .A(n11257), .B(U157_Z_2), .Z(n11256) );
  AN2 U7416 ( .A(n11105), .B(n11258), .Z(n11255) );
  OR2 U7417 ( .A(n11108), .B(n11128), .Z(n11258) );
  OR2 U7418 ( .A(n8835), .B(n8831), .Z(n11128) );
  AN2 U7419 ( .A(n11259), .B(n11260), .Z(n8831) );
  AN2 U7420 ( .A(n5329), .B(n1704), .Z(n11260) );
  IV U7421 ( .A(n1648), .Z(n5329) );
  AN2 U7422 ( .A(n5330), .B(n11179), .Z(n8835) );
  AN2 U7423 ( .A(n11259), .B(n11261), .Z(n11179) );
  AN2 U7424 ( .A(n1648), .B(n1704), .Z(n11261) );
  IV U7425 ( .A(n1596), .Z(n5330) );
  OR2 U7426 ( .A(n8834), .B(n8832), .Z(n11108) );
  AN2 U7427 ( .A(n5328), .B(n11259), .Z(n8832) );
  AN2 U7428 ( .A(U154_Z_0), .B(n11262), .Z(n11259) );
  AN2 U7429 ( .A(n1768), .B(n1809), .Z(n11262) );
  IV U7430 ( .A(n1704), .Z(n5328) );
  AN2 U7431 ( .A(U154_Z_0), .B(n11263), .Z(n8834) );
  AN2 U7432 ( .A(n5327), .B(n1809), .Z(n11263) );
  IV U7433 ( .A(n1768), .Z(n5327) );
  AN2 U7434 ( .A(n10125), .B(n11086), .Z(n11105) );
  OR2 U7435 ( .A(n8731), .B(n11264), .Z(n11086) );
  AN2 U7436 ( .A(n10856), .B(U156_Z_6), .Z(n11253) );
  OR2 U7437 ( .A(n11265), .B(n11266), .Z(tx_data_out[16]) );
  AN2 U7438 ( .A(n9942), .B(n11267), .Z(n11266) );
  AN2 U7439 ( .A(n9929), .B(n9212), .Z(n11265) );
  OR2 U7440 ( .A(n11268), .B(n11269), .Z(n9212) );
  AN2 U7441 ( .A(n11270), .B(n11271), .Z(n11269) );
  IV U7442 ( .A(U37_DATA1_14), .Z(n11271) );
  AN2 U7443 ( .A(n11272), .B(U37_DATA1_14), .Z(n11268) );
  IV U7444 ( .A(n11270), .Z(n11272) );
  OR2 U7445 ( .A(n11273), .B(n11274), .Z(n11270) );
  AN2 U7446 ( .A(n11275), .B(n10787), .Z(n11274) );
  IV U7447 ( .A(U37_DATA1_33), .Z(n10787) );
  OR2 U7448 ( .A(n11276), .B(n1934), .Z(n11275) );
  AN2 U7449 ( .A(n11267), .B(n5684), .Z(n11276) );
  AN2 U7450 ( .A(U37_DATA1_33), .B(n11277), .Z(n11273) );
  OR2 U7451 ( .A(n11278), .B(n9953), .Z(n11277) );
  AN2 U7452 ( .A(n11279), .B(n9955), .Z(n11278) );
  IV U7453 ( .A(n11267), .Z(n11279) );
  OR2 U7454 ( .A(n11280), .B(n11281), .Z(n11267) );
  OR2 U7455 ( .A(n11282), .B(n11283), .Z(n11281) );
  AN2 U7456 ( .A(n11257), .B(U156_Z_1), .Z(n11283) );
  AN2 U7457 ( .A(n11284), .B(n11285), .Z(n11282) );
  OR2 U7458 ( .A(n8846), .B(n11286), .Z(n11285) );
  OR2 U7459 ( .A(n8843), .B(n11287), .Z(n11286) );
  AN2 U7460 ( .A(n10856), .B(U156_Z_5), .Z(n11280) );
  OR2 U7461 ( .A(n11288), .B(n11289), .Z(tx_data_out[15]) );
  AN2 U7462 ( .A(n9942), .B(n11290), .Z(n11289) );
  AN2 U7463 ( .A(n9929), .B(n9223), .Z(n11288) );
  OR2 U7464 ( .A(n11291), .B(n11292), .Z(n9223) );
  AN2 U7465 ( .A(n11293), .B(n11294), .Z(n11292) );
  IV U7466 ( .A(U37_DATA1_13), .Z(n11294) );
  AN2 U7467 ( .A(n11295), .B(U37_DATA1_13), .Z(n11291) );
  IV U7468 ( .A(n11293), .Z(n11295) );
  OR2 U7469 ( .A(n11296), .B(n11297), .Z(n11293) );
  AN2 U7470 ( .A(n11298), .B(n10814), .Z(n11297) );
  IV U7471 ( .A(U37_DATA1_32), .Z(n10814) );
  OR2 U7472 ( .A(n11299), .B(n1934), .Z(n11298) );
  AN2 U7473 ( .A(n11290), .B(n5684), .Z(n11299) );
  AN2 U7474 ( .A(U37_DATA1_32), .B(n11300), .Z(n11296) );
  OR2 U7475 ( .A(n11301), .B(n9953), .Z(n11300) );
  AN2 U7476 ( .A(n11302), .B(n9955), .Z(n11301) );
  IV U7477 ( .A(n11290), .Z(n11302) );
  OR2 U7478 ( .A(n11303), .B(n11304), .Z(n11290) );
  OR2 U7479 ( .A(n11305), .B(n11306), .Z(n11304) );
  AN2 U7480 ( .A(n11257), .B(U156_Z_0), .Z(n11306) );
  AN2 U7481 ( .A(n11284), .B(n11307), .Z(n11305) );
  OR2 U7482 ( .A(n8847), .B(n11308), .Z(n11307) );
  OR2 U7483 ( .A(n8844), .B(n11287), .Z(n11308) );
  AN2 U7484 ( .A(n11309), .B(n8850), .Z(n11287) );
  AN2 U7485 ( .A(n10856), .B(U156_Z_4), .Z(n11303) );
  OR2 U7486 ( .A(n11310), .B(n11311), .Z(tx_data_out[14]) );
  OR2 U7487 ( .A(n11312), .B(n11313), .Z(n11311) );
  AN2 U7488 ( .A(n9930), .B(n11314), .Z(n11313) );
  AN2 U7489 ( .A(n9929), .B(n9234), .Z(n11312) );
  AN2 U7490 ( .A(n11315), .B(n11316), .Z(n9234) );
  IV U7491 ( .A(n11317), .Z(n11316) );
  AN2 U7492 ( .A(n11318), .B(n11319), .Z(n11317) );
  OR2 U7493 ( .A(n11319), .B(n11318), .Z(n11315) );
  OR2 U7494 ( .A(n11320), .B(n11321), .Z(n11318) );
  AN2 U7495 ( .A(U37_DATA1_12), .B(n10843), .Z(n11321) );
  IV U7496 ( .A(U37_DATA1_31), .Z(n10843) );
  AN2 U7497 ( .A(U37_DATA1_31), .B(n11322), .Z(n11320) );
  IV U7498 ( .A(U37_DATA1_12), .Z(n11322) );
  OR2 U7499 ( .A(n11323), .B(n11324), .Z(n11319) );
  OR2 U7500 ( .A(n1934), .B(n11325), .Z(n11324) );
  AN2 U7501 ( .A(n10414), .B(n11314), .Z(n11325) );
  OR2 U7502 ( .A(n11326), .B(n11327), .Z(n11314) );
  OR2 U7503 ( .A(n11328), .B(n11329), .Z(n11327) );
  AN2 U7504 ( .A(n1907), .B(U157_Z_1), .Z(n11328) );
  OR2 U7505 ( .A(n11330), .B(n11331), .Z(n11326) );
  AN2 U7506 ( .A(n8735), .B(U156_Z_3), .Z(n11331) );
  AN2 U7507 ( .A(n11332), .B(n11264), .Z(n11330) );
  AN2 U7508 ( .A(n10413), .B(U156_Z_3), .Z(n11323) );
  AN2 U7509 ( .A(n9928), .B(U156_Z_3), .Z(n11310) );
  OR2 U7510 ( .A(n11333), .B(n11334), .Z(tx_data_out[13]) );
  OR2 U7511 ( .A(n11335), .B(n11336), .Z(n11334) );
  AN2 U7512 ( .A(n9930), .B(n11337), .Z(n11336) );
  AN2 U7513 ( .A(n9929), .B(n9333), .Z(n11335) );
  AN2 U7514 ( .A(n11338), .B(n11339), .Z(n9333) );
  IV U7515 ( .A(n11340), .Z(n11339) );
  AN2 U7516 ( .A(n11341), .B(n11342), .Z(n11340) );
  OR2 U7517 ( .A(n11342), .B(n11341), .Z(n11338) );
  OR2 U7518 ( .A(n11343), .B(n11344), .Z(n11341) );
  AN2 U7519 ( .A(U37_DATA1_11), .B(n10865), .Z(n11344) );
  IV U7520 ( .A(U37_DATA1_30), .Z(n10865) );
  AN2 U7521 ( .A(U37_DATA1_30), .B(n11345), .Z(n11343) );
  IV U7522 ( .A(U37_DATA1_11), .Z(n11345) );
  OR2 U7523 ( .A(n11346), .B(n11347), .Z(n11342) );
  OR2 U7524 ( .A(n1934), .B(n11348), .Z(n11347) );
  AN2 U7525 ( .A(n10413), .B(U156_Z_2), .Z(n11348) );
  AN2 U7526 ( .A(n5684), .B(n99), .Z(n10413) );
  AN2 U7527 ( .A(n10414), .B(n11337), .Z(n11346) );
  OR2 U7528 ( .A(n11349), .B(n11350), .Z(n11337) );
  OR2 U7529 ( .A(n11351), .B(n11329), .Z(n11350) );
  OR2 U7530 ( .A(n11352), .B(n8755), .Z(n11329) );
  AN2 U7531 ( .A(n11353), .B(n11264), .Z(n11352) );
  OR2 U7532 ( .A(n11354), .B(n11355), .Z(n11353) );
  AN2 U7533 ( .A(n8851), .B(n11356), .Z(n11355) );
  OR2 U7534 ( .A(n1327), .B(n5313), .Z(n11356) );
  IV U7535 ( .A(n1433), .Z(n5313) );
  AN2 U7536 ( .A(n11357), .B(n8850), .Z(n8851) );
  IV U7537 ( .A(n11309), .Z(n11357) );
  OR2 U7538 ( .A(n5312), .B(n5305), .Z(n11309) );
  IV U7539 ( .A(n1554), .Z(n5312) );
  AN2 U7540 ( .A(n11358), .B(n8850), .Z(n11354) );
  AN2 U7541 ( .A(n1610), .B(n11359), .Z(n8850) );
  AN2 U7542 ( .A(n1554), .B(n5305), .Z(n11358) );
  IV U7543 ( .A(n1492), .Z(n5305) );
  AN2 U7544 ( .A(n1907), .B(U157_Z_0), .Z(n11351) );
  OR2 U7545 ( .A(n11360), .B(n11361), .Z(n11349) );
  AN2 U7546 ( .A(n8735), .B(U156_Z_2), .Z(n11361) );
  AN2 U7547 ( .A(n11362), .B(n11264), .Z(n11360) );
  AN2 U7548 ( .A(n10125), .B(n5684), .Z(n10414) );
  AN2 U7549 ( .A(n9928), .B(U156_Z_2), .Z(n11333) );
  OR2 U7550 ( .A(n11363), .B(n11364), .Z(tx_data_out[12]) );
  AN2 U7551 ( .A(n9942), .B(n11365), .Z(n11364) );
  AN2 U7552 ( .A(n9929), .B(n9454), .Z(n11363) );
  OR2 U7553 ( .A(n11366), .B(n11367), .Z(n9454) );
  AN2 U7554 ( .A(n11368), .B(n11369), .Z(n11367) );
  IV U7555 ( .A(U37_DATA1_10), .Z(n11369) );
  AN2 U7556 ( .A(n11370), .B(U37_DATA1_10), .Z(n11366) );
  IV U7557 ( .A(n11368), .Z(n11370) );
  OR2 U7558 ( .A(n11371), .B(n11372), .Z(n11368) );
  AN2 U7559 ( .A(n11373), .B(n10885), .Z(n11372) );
  IV U7560 ( .A(U37_DATA1_29), .Z(n10885) );
  OR2 U7561 ( .A(n11374), .B(n1934), .Z(n11373) );
  AN2 U7562 ( .A(n11365), .B(n5684), .Z(n11374) );
  AN2 U7563 ( .A(U37_DATA1_29), .B(n11375), .Z(n11371) );
  OR2 U7564 ( .A(n11376), .B(n9953), .Z(n11375) );
  AN2 U7565 ( .A(n11377), .B(n9955), .Z(n11376) );
  IV U7566 ( .A(n11365), .Z(n11377) );
  OR2 U7567 ( .A(n11378), .B(n11379), .Z(n11365) );
  OR2 U7568 ( .A(n11380), .B(n11381), .Z(n11379) );
  AN2 U7569 ( .A(U59_DATA1_1), .B(n11284), .Z(n11381) );
  AN2 U7570 ( .A(n11257), .B(U159_Z_1), .Z(n11380) );
  OR2 U7571 ( .A(n10038), .B(n11382), .Z(n11378) );
  AN2 U7572 ( .A(n10856), .B(n8672), .Z(n11382) );
  OR2 U7573 ( .A(n11383), .B(n4170), .Z(n8672) );
  AN2 U7574 ( .A(U162_DATA3_10), .B(n10092), .Z(n11383) );
  OR2 U7575 ( .A(n11384), .B(n11385), .Z(tx_data_out[11]) );
  AN2 U7576 ( .A(n9942), .B(n11386), .Z(n11385) );
  AN2 U7577 ( .A(n9929), .B(n9575), .Z(n11384) );
  OR2 U7578 ( .A(n11387), .B(n11388), .Z(n9575) );
  AN2 U7579 ( .A(n11389), .B(n11390), .Z(n11388) );
  IV U7580 ( .A(U37_DATA1_9), .Z(n11390) );
  AN2 U7581 ( .A(n11391), .B(U37_DATA1_9), .Z(n11387) );
  IV U7582 ( .A(n11389), .Z(n11391) );
  OR2 U7583 ( .A(n11392), .B(n11393), .Z(n11389) );
  AN2 U7584 ( .A(n11394), .B(n10910), .Z(n11393) );
  IV U7585 ( .A(U37_DATA1_28), .Z(n10910) );
  OR2 U7586 ( .A(n11395), .B(n1934), .Z(n11394) );
  AN2 U7587 ( .A(n11386), .B(n5684), .Z(n11395) );
  AN2 U7588 ( .A(U37_DATA1_28), .B(n11396), .Z(n11392) );
  OR2 U7589 ( .A(n11397), .B(n9953), .Z(n11396) );
  AN2 U7590 ( .A(n11398), .B(n9955), .Z(n11397) );
  IV U7591 ( .A(n11386), .Z(n11398) );
  OR2 U7592 ( .A(n11399), .B(n11400), .Z(n11386) );
  OR2 U7593 ( .A(n11401), .B(n11402), .Z(n11400) );
  AN2 U7594 ( .A(n10856), .B(U158_Z_1), .Z(n11402) );
  AN2 U7595 ( .A(U59_DATA1_0), .B(n11284), .Z(n11401) );
  OR2 U7596 ( .A(n10038), .B(n11403), .Z(n11399) );
  AN2 U7597 ( .A(n11257), .B(U158_Z_0), .Z(n11403) );
  AN2 U7598 ( .A(n10125), .B(n8755), .Z(n10038) );
  IV U7599 ( .A(n11404), .Z(n8755) );
  OR2 U7600 ( .A(n11405), .B(n11406), .Z(n11404) );
  OR2 U7601 ( .A(n8737), .B(n10986), .Z(n11406) );
  OR2 U7602 ( .A(n8728), .B(n10771), .Z(n10986) );
  OR2 U7603 ( .A(n1929), .B(n5245), .Z(n10771) );
  IV U7604 ( .A(n11407), .Z(n5245) );
  OR2 U7605 ( .A(n643), .B(n644), .Z(n11407) );
  OR2 U7606 ( .A(n5247), .B(n11408), .Z(n1929) );
  OR2 U7607 ( .A(n5246), .B(n5248), .Z(n11408) );
  IV U7608 ( .A(n11409), .Z(n5248) );
  OR2 U7609 ( .A(n595), .B(n596), .Z(n11409) );
  IV U7610 ( .A(n11410), .Z(n5246) );
  OR2 U7611 ( .A(n628), .B(n627), .Z(n11410) );
  IV U7612 ( .A(n11411), .Z(n5247) );
  OR2 U7613 ( .A(n611), .B(n612), .Z(n11411) );
  IV U7614 ( .A(n11412), .Z(n8728) );
  OR2 U7615 ( .A(n579), .B(n580), .Z(n11412) );
  OR2 U7616 ( .A(n8758), .B(n11413), .Z(n8737) );
  OR2 U7617 ( .A(n8753), .B(n8742), .Z(n11413) );
  OR2 U7618 ( .A(n1918), .B(n5254), .Z(n11405) );
  OR2 U7619 ( .A(n11414), .B(n8757), .Z(n1918) );
  OR2 U7620 ( .A(n8731), .B(n8748), .Z(n8757) );
  OR2 U7621 ( .A(n11415), .B(n8744), .Z(n8748) );
  IV U7622 ( .A(n11416), .Z(n8731) );
  OR2 U7623 ( .A(n531), .B(n532), .Z(n11416) );
  OR2 U7624 ( .A(n5249), .B(n8734), .Z(n11414) );
  IV U7625 ( .A(n11417), .Z(n8734) );
  OR2 U7626 ( .A(n547), .B(n548), .Z(n11417) );
  IV U7627 ( .A(n11418), .Z(n5249) );
  OR2 U7628 ( .A(n563), .B(n564), .Z(n11418) );
  OR2 U7629 ( .A(n11419), .B(n11420), .Z(tx_data_out[10]) );
  AN2 U7630 ( .A(n9942), .B(n11421), .Z(n11420) );
  AN2 U7631 ( .A(n9929), .B(n9696), .Z(n11419) );
  OR2 U7632 ( .A(n11422), .B(n11423), .Z(n9696) );
  AN2 U7633 ( .A(n11424), .B(n11425), .Z(n11423) );
  IV U7634 ( .A(U37_DATA1_8), .Z(n11425) );
  AN2 U7635 ( .A(n11426), .B(U37_DATA1_8), .Z(n11422) );
  IV U7636 ( .A(n11424), .Z(n11426) );
  OR2 U7637 ( .A(n11427), .B(n11428), .Z(n11424) );
  AN2 U7638 ( .A(n11429), .B(n10949), .Z(n11428) );
  IV U7639 ( .A(U37_DATA1_27), .Z(n10949) );
  OR2 U7640 ( .A(n11430), .B(n1934), .Z(n11429) );
  AN2 U7641 ( .A(n11421), .B(n5684), .Z(n11430) );
  IV U7642 ( .A(n98), .Z(n5684) );
  AN2 U7643 ( .A(U37_DATA1_27), .B(n11431), .Z(n11427) );
  OR2 U7644 ( .A(n11432), .B(n9953), .Z(n11431) );
  AN2 U7645 ( .A(n9955), .B(n98), .Z(n9953) );
  AN2 U7646 ( .A(n11433), .B(n9955), .Z(n11432) );
  IV U7647 ( .A(n1934), .Z(n9955) );
  IV U7648 ( .A(n11421), .Z(n11433) );
  OR2 U7649 ( .A(n11434), .B(n11435), .Z(n11421) );
  OR2 U7650 ( .A(n11436), .B(n11437), .Z(n11435) );
  AN2 U7651 ( .A(n11257), .B(U159_Z_0), .Z(n11437) );
  AN2 U7652 ( .A(n10125), .B(n1907), .Z(n11257) );
  AN2 U7653 ( .A(n11284), .B(n11438), .Z(n11436) );
  OR2 U7654 ( .A(n11362), .B(n11332), .Z(n11438) );
  OR2 U7655 ( .A(n8847), .B(n8843), .Z(n11332) );
  AN2 U7656 ( .A(n5309), .B(n11439), .Z(n8843) );
  IV U7657 ( .A(n1720), .Z(n5309) );
  AN2 U7658 ( .A(n5311), .B(n11359), .Z(n8847) );
  AN2 U7659 ( .A(n11439), .B(n11440), .Z(n11359) );
  AN2 U7660 ( .A(n1660), .B(n1720), .Z(n11440) );
  IV U7661 ( .A(n1610), .Z(n5311) );
  OR2 U7662 ( .A(n8846), .B(n8844), .Z(n11362) );
  AN2 U7663 ( .A(n11439), .B(n11441), .Z(n8844) );
  AN2 U7664 ( .A(n5310), .B(n1720), .Z(n11441) );
  IV U7665 ( .A(n1660), .Z(n5310) );
  AN2 U7666 ( .A(U155_Z_0), .B(n11442), .Z(n11439) );
  AN2 U7667 ( .A(n1783), .B(n1815), .Z(n11442) );
  AN2 U7668 ( .A(U155_Z_0), .B(n11443), .Z(n8846) );
  AN2 U7669 ( .A(n5308), .B(n1815), .Z(n11443) );
  IV U7670 ( .A(n1783), .Z(n5308) );
  AN2 U7671 ( .A(n10125), .B(n11264), .Z(n11284) );
  OR2 U7672 ( .A(n8744), .B(n8758), .Z(n11264) );
  OR2 U7673 ( .A(n8745), .B(n5257), .Z(n8758) );
  IV U7674 ( .A(n11444), .Z(n5257) );
  OR2 U7675 ( .A(n436), .B(n435), .Z(n11444) );
  IV U7676 ( .A(n11445), .Z(n8745) );
  OR2 U7677 ( .A(n452), .B(n451), .Z(n11445) );
  IV U7678 ( .A(n11446), .Z(n8744) );
  OR2 U7679 ( .A(n420), .B(n419), .Z(n11446) );
  AN2 U7680 ( .A(n10856), .B(U159_Z_2), .Z(n11434) );
  OR2 U7681 ( .A(n99), .B(n8735), .Z(n10856) );
  OR2 U7682 ( .A(n8742), .B(n10767), .Z(n8735) );
  OR2 U7683 ( .A(n8753), .B(n8760), .Z(n10767) );
  OR2 U7684 ( .A(n11415), .B(n5254), .Z(n8760) );
  IV U7685 ( .A(n11447), .Z(n5254) );
  OR2 U7686 ( .A(n483), .B(n484), .Z(n11447) );
  AN2 U7687 ( .A(n11448), .B(n11449), .Z(n11415) );
  IV U7688 ( .A(n516), .Z(n11449) );
  IV U7689 ( .A(n515), .Z(n11448) );
  IV U7690 ( .A(n11450), .Z(n8753) );
  OR2 U7691 ( .A(n468), .B(n467), .Z(n11450) );
  IV U7692 ( .A(n11451), .Z(n8742) );
  OR2 U7693 ( .A(n499), .B(n500), .Z(n11451) );
  OR2 U7694 ( .A(n11452), .B(n9928), .Z(tx_data_out[1]) );
  AN2 U7695 ( .A(n99), .B(n9942), .Z(n9928) );
  AN2 U7696 ( .A(n9929), .B(n99), .Z(n11452) );
  OR2 U7697 ( .A(n11453), .B(n9930), .Z(tx_data_out[0]) );
  AN2 U7698 ( .A(n10125), .B(n9942), .Z(n9930) );
  AN2 U7699 ( .A(U107_DATA1_0), .B(n11454), .Z(n9942) );
  IV U7700 ( .A(n11455), .Z(n11454) );
  AN2 U7701 ( .A(n9929), .B(n10125), .Z(n11453) );
  IV U7702 ( .A(n99), .Z(n10125) );
  IV U7703 ( .A(n11456), .Z(n9929) );
  OR2 U7704 ( .A(U107_DATA1_0), .B(n11455), .Z(n11456) );
  OR2 U7705 ( .A(n4614), .B(n4479), .Z(n11455) );
  OR2 U7706 ( .A(n11457), .B(n8179), .Z(U162_Z_9) );
  AN2 U7707 ( .A(U161_CONTROL3), .B(U162_DATA3_9), .Z(n11457) );
  OR2 U7708 ( .A(n11458), .B(n8182), .Z(U162_Z_8) );
  AN2 U7709 ( .A(U161_CONTROL3), .B(U162_DATA3_8), .Z(n11458) );
  OR2 U7710 ( .A(n11459), .B(n8184), .Z(U162_Z_7) );
  AN2 U7711 ( .A(U161_CONTROL3), .B(U162_DATA3_7), .Z(n11459) );
  OR2 U7712 ( .A(n11460), .B(n8186), .Z(U162_Z_63) );
  AN2 U7713 ( .A(U161_CONTROL3), .B(U162_DATA3_63), .Z(n11460) );
  OR2 U7714 ( .A(n11461), .B(n8188), .Z(U162_Z_62) );
  AN2 U7715 ( .A(U161_CONTROL3), .B(U162_DATA3_62), .Z(n11461) );
  OR2 U7716 ( .A(n11462), .B(n8190), .Z(U162_Z_61) );
  AN2 U7717 ( .A(U161_CONTROL3), .B(U162_DATA3_61), .Z(n11462) );
  OR2 U7718 ( .A(n11463), .B(n8192), .Z(U162_Z_60) );
  AN2 U7719 ( .A(U161_CONTROL3), .B(U162_DATA3_60), .Z(n11463) );
  OR2 U7720 ( .A(n11464), .B(n8194), .Z(U162_Z_6) );
  AN2 U7721 ( .A(U161_CONTROL3), .B(U162_DATA3_6), .Z(n11464) );
  OR2 U7722 ( .A(n11465), .B(n8196), .Z(U162_Z_59) );
  AN2 U7723 ( .A(U161_CONTROL3), .B(U162_DATA3_59), .Z(n11465) );
  OR2 U7724 ( .A(n11466), .B(n8199), .Z(U162_Z_58) );
  AN2 U7725 ( .A(U161_CONTROL3), .B(U162_DATA3_58), .Z(n11466) );
  OR2 U7726 ( .A(n11467), .B(n8202), .Z(U162_Z_57) );
  AN2 U7727 ( .A(U161_CONTROL3), .B(U162_DATA3_57), .Z(n11467) );
  OR2 U7728 ( .A(n11468), .B(n8205), .Z(U162_Z_56) );
  AN2 U7729 ( .A(U161_CONTROL3), .B(U162_DATA3_56), .Z(n11468) );
  OR2 U7730 ( .A(n11469), .B(n8207), .Z(U162_Z_55) );
  AN2 U7731 ( .A(U161_CONTROL3), .B(U162_DATA3_55), .Z(n11469) );
  OR2 U7732 ( .A(n11470), .B(n8209), .Z(U162_Z_54) );
  AN2 U7733 ( .A(U161_CONTROL3), .B(U162_DATA3_54), .Z(n11470) );
  OR2 U7734 ( .A(n11471), .B(n8211), .Z(U162_Z_53) );
  AN2 U7735 ( .A(U161_CONTROL3), .B(U162_DATA3_53), .Z(n11471) );
  OR2 U7736 ( .A(n11472), .B(n8213), .Z(U162_Z_52) );
  AN2 U7737 ( .A(U161_CONTROL3), .B(U162_DATA3_52), .Z(n11472) );
  OR2 U7738 ( .A(n11473), .B(n8215), .Z(U162_Z_51) );
  AN2 U7739 ( .A(U161_CONTROL3), .B(U162_DATA3_51), .Z(n11473) );
  OR2 U7740 ( .A(n11474), .B(n8218), .Z(U162_Z_50) );
  AN2 U7741 ( .A(U161_CONTROL3), .B(U162_DATA3_50), .Z(n11474) );
  OR2 U7742 ( .A(n11475), .B(n8220), .Z(U162_Z_5) );
  AN2 U7743 ( .A(U161_CONTROL3), .B(U162_DATA3_5), .Z(n11475) );
  OR2 U7744 ( .A(n11476), .B(n8223), .Z(U162_Z_49) );
  AN2 U7745 ( .A(U161_CONTROL3), .B(U162_DATA3_49), .Z(n11476) );
  OR2 U7746 ( .A(n11477), .B(n8226), .Z(U162_Z_48) );
  AN2 U7747 ( .A(U161_CONTROL3), .B(U162_DATA3_48), .Z(n11477) );
  OR2 U7748 ( .A(n11478), .B(n8228), .Z(U162_Z_47) );
  AN2 U7749 ( .A(U161_CONTROL3), .B(U162_DATA3_47), .Z(n11478) );
  OR2 U7750 ( .A(n11479), .B(n8230), .Z(U162_Z_46) );
  AN2 U7751 ( .A(U161_CONTROL3), .B(U162_DATA3_46), .Z(n11479) );
  OR2 U7752 ( .A(n11480), .B(n8232), .Z(U162_Z_45) );
  AN2 U7753 ( .A(U161_CONTROL3), .B(U162_DATA3_45), .Z(n11480) );
  OR2 U7754 ( .A(n11481), .B(n8234), .Z(U162_Z_44) );
  AN2 U7755 ( .A(U161_CONTROL3), .B(U162_DATA3_44), .Z(n11481) );
  OR2 U7756 ( .A(n11482), .B(n8236), .Z(U162_Z_43) );
  AN2 U7757 ( .A(U161_CONTROL3), .B(U162_DATA3_43), .Z(n11482) );
  OR2 U7758 ( .A(n11483), .B(n8239), .Z(U162_Z_42) );
  AN2 U7759 ( .A(U161_CONTROL3), .B(U162_DATA3_42), .Z(n11483) );
  OR2 U7760 ( .A(n11484), .B(n8242), .Z(U162_Z_41) );
  AN2 U7761 ( .A(U161_CONTROL3), .B(U162_DATA3_41), .Z(n11484) );
  OR2 U7762 ( .A(n11485), .B(n8245), .Z(U162_Z_40) );
  AN2 U7763 ( .A(U161_CONTROL3), .B(U162_DATA3_40), .Z(n11485) );
  OR2 U7764 ( .A(n11486), .B(n8247), .Z(U162_Z_4) );
  AN2 U7765 ( .A(U161_CONTROL3), .B(U162_DATA3_4), .Z(n11486) );
  OR2 U7766 ( .A(n11487), .B(n8249), .Z(U162_Z_39) );
  AN2 U7767 ( .A(U161_CONTROL3), .B(U162_DATA3_39), .Z(n11487) );
  OR2 U7768 ( .A(n11488), .B(n8251), .Z(U162_Z_38) );
  AN2 U7769 ( .A(U161_CONTROL3), .B(U162_DATA3_38), .Z(n11488) );
  OR2 U7770 ( .A(n11489), .B(n8253), .Z(U162_Z_37) );
  AN2 U7771 ( .A(U161_CONTROL3), .B(U162_DATA3_37), .Z(n11489) );
  OR2 U7772 ( .A(n11490), .B(n8255), .Z(U162_Z_36) );
  AN2 U7773 ( .A(U161_CONTROL3), .B(U162_DATA3_36), .Z(n11490) );
  OR2 U7774 ( .A(n11491), .B(n8257), .Z(U162_Z_35) );
  AN2 U7775 ( .A(U161_CONTROL3), .B(U162_DATA3_35), .Z(n11491) );
  OR2 U7776 ( .A(n11492), .B(n8260), .Z(U162_Z_34) );
  AN2 U7777 ( .A(U162_DATA3_34), .B(U161_CONTROL3), .Z(n11492) );
  OR2 U7778 ( .A(n11493), .B(n8263), .Z(U162_Z_33) );
  AN2 U7779 ( .A(U161_CONTROL3), .B(U162_DATA3_33), .Z(n11493) );
  OR2 U7780 ( .A(n11494), .B(n8266), .Z(U162_Z_32) );
  AN2 U7781 ( .A(U161_CONTROL3), .B(U162_DATA3_32), .Z(n11494) );
  OR2 U7782 ( .A(n11495), .B(n8268), .Z(U162_Z_31) );
  AN2 U7783 ( .A(U161_CONTROL3), .B(U162_DATA3_31), .Z(n11495) );
  OR2 U7784 ( .A(n11496), .B(n8270), .Z(U162_Z_30) );
  AN2 U7785 ( .A(U161_CONTROL3), .B(U162_DATA3_30), .Z(n11496) );
  OR2 U7786 ( .A(n11497), .B(n8272), .Z(U162_Z_3) );
  AN2 U7787 ( .A(U161_CONTROL3), .B(U162_DATA3_3), .Z(n11497) );
  OR2 U7788 ( .A(n11498), .B(n8274), .Z(U162_Z_29) );
  AN2 U7789 ( .A(U161_CONTROL3), .B(U162_DATA3_29), .Z(n11498) );
  OR2 U7790 ( .A(n11499), .B(n8276), .Z(U162_Z_28) );
  AN2 U7791 ( .A(U161_CONTROL3), .B(U162_DATA3_28), .Z(n11499) );
  OR2 U7792 ( .A(n11500), .B(n8278), .Z(U162_Z_27) );
  AN2 U7793 ( .A(U161_CONTROL3), .B(U162_DATA3_27), .Z(n11500) );
  OR2 U7794 ( .A(n11501), .B(n8281), .Z(U162_Z_26) );
  AN2 U7795 ( .A(U161_CONTROL3), .B(U162_DATA3_26), .Z(n11501) );
  OR2 U7796 ( .A(n11502), .B(n8284), .Z(U162_Z_25) );
  AN2 U7797 ( .A(U161_CONTROL3), .B(U162_DATA3_25), .Z(n11502) );
  OR2 U7798 ( .A(n11503), .B(n8287), .Z(U162_Z_24) );
  AN2 U7799 ( .A(U161_CONTROL3), .B(U162_DATA3_24), .Z(n11503) );
  OR2 U7800 ( .A(n11504), .B(n8289), .Z(U162_Z_23) );
  AN2 U7801 ( .A(U161_CONTROL3), .B(U162_DATA3_23), .Z(n11504) );
  OR2 U7802 ( .A(n11505), .B(n8291), .Z(U162_Z_22) );
  AN2 U7803 ( .A(U161_CONTROL3), .B(U162_DATA3_22), .Z(n11505) );
  OR2 U7804 ( .A(n11506), .B(n8293), .Z(U162_Z_21) );
  AN2 U7805 ( .A(U161_CONTROL3), .B(U162_DATA3_21), .Z(n11506) );
  OR2 U7806 ( .A(n11507), .B(n8295), .Z(U162_Z_20) );
  AN2 U7807 ( .A(U161_CONTROL3), .B(U162_DATA3_20), .Z(n11507) );
  OR2 U7808 ( .A(n11508), .B(n8298), .Z(U162_Z_2) );
  AN2 U7809 ( .A(U162_DATA3_2), .B(U161_CONTROL3), .Z(n11508) );
  OR2 U7810 ( .A(n11509), .B(n8300), .Z(U162_Z_19) );
  AN2 U7811 ( .A(U161_CONTROL3), .B(U162_DATA3_19), .Z(n11509) );
  OR2 U7812 ( .A(n11510), .B(n8303), .Z(U162_Z_18) );
  AN2 U7813 ( .A(U161_CONTROL3), .B(U162_DATA3_18), .Z(n11510) );
  OR2 U7814 ( .A(n11511), .B(n8306), .Z(U162_Z_17) );
  AN2 U7815 ( .A(U161_CONTROL3), .B(U162_DATA3_17), .Z(n11511) );
  OR2 U7816 ( .A(n11512), .B(n8309), .Z(U162_Z_16) );
  AN2 U7817 ( .A(U161_CONTROL3), .B(U162_DATA3_16), .Z(n11512) );
  OR2 U7818 ( .A(n11513), .B(n8311), .Z(U162_Z_15) );
  AN2 U7819 ( .A(U161_CONTROL3), .B(U162_DATA3_15), .Z(n11513) );
  OR2 U7820 ( .A(n11514), .B(n8313), .Z(U162_Z_14) );
  AN2 U7821 ( .A(U161_CONTROL3), .B(U162_DATA3_14), .Z(n11514) );
  OR2 U7822 ( .A(n11515), .B(n8315), .Z(U162_Z_13) );
  AN2 U7823 ( .A(U161_CONTROL3), .B(U162_DATA3_13), .Z(n11515) );
  OR2 U7824 ( .A(n11516), .B(n8317), .Z(U162_Z_12) );
  AN2 U7825 ( .A(U161_CONTROL3), .B(U162_DATA3_12), .Z(n11516) );
  OR2 U7826 ( .A(n11517), .B(n8319), .Z(U162_Z_11) );
  AN2 U7827 ( .A(U161_CONTROL3), .B(U162_DATA3_11), .Z(n11517) );
  OR2 U7828 ( .A(n11518), .B(n8322), .Z(U162_Z_10) );
  AN2 U7829 ( .A(U161_CONTROL3), .B(U162_DATA3_10), .Z(n11518) );
  OR2 U7830 ( .A(n11519), .B(n8325), .Z(U162_Z_1) );
  AN2 U7831 ( .A(U161_CONTROL3), .B(U162_DATA3_1), .Z(n11519) );
  OR2 U7832 ( .A(n11520), .B(n8328), .Z(U162_Z_0) );
  AN2 U7833 ( .A(U161_CONTROL3), .B(U162_DATA3_0), .Z(n11520) );
  OR2 U7834 ( .A(n11521), .B(n8331), .Z(U161_Z_7) );
  AN2 U7835 ( .A(U161_CONTROL3), .B(U161_DATA3_7), .Z(n11521) );
  OR2 U7836 ( .A(n11522), .B(n8334), .Z(U161_Z_6) );
  AN2 U7837 ( .A(U161_CONTROL3), .B(U161_DATA3_6), .Z(n11522) );
  OR2 U7838 ( .A(n11523), .B(n8337), .Z(U161_Z_5) );
  AN2 U7839 ( .A(U161_CONTROL3), .B(U161_DATA3_5), .Z(n11523) );
  OR2 U7840 ( .A(n11524), .B(n8340), .Z(U161_Z_4) );
  AN2 U7841 ( .A(U161_DATA3_4), .B(U161_CONTROL3), .Z(n11524) );
  OR2 U7842 ( .A(n11525), .B(n8343), .Z(U161_Z_3) );
  AN2 U7843 ( .A(U161_CONTROL3), .B(U161_DATA3_3), .Z(n11525) );
  OR2 U7844 ( .A(n11526), .B(n8346), .Z(U161_Z_2) );
  AN2 U7845 ( .A(U161_CONTROL3), .B(U161_DATA3_2), .Z(n11526) );
  OR2 U7846 ( .A(n11527), .B(n8349), .Z(U161_Z_1) );
  AN2 U7847 ( .A(U161_CONTROL3), .B(U161_DATA3_1), .Z(n11527) );
  OR2 U7848 ( .A(n11528), .B(n8352), .Z(U161_Z_0) );
  AN2 U7849 ( .A(U161_DATA3_0), .B(U161_CONTROL3), .Z(n11528) );
  OR2 U7850 ( .A(n11529), .B(reset_to_pma_tx), .Z(U160_Z_3) );
  AN2 U7851 ( .A(n3179), .B(U160_DATA2_3), .Z(n11529) );
  OR2 U7852 ( .A(n11530), .B(reset_to_pma_tx), .Z(U160_Z_2) );
  AN2 U7853 ( .A(n3179), .B(U160_DATA2_2), .Z(n11530) );
  OR2 U7854 ( .A(n11531), .B(reset_to_pma_tx), .Z(U160_Z_1) );
  AN2 U7855 ( .A(n3179), .B(U160_DATA2_1), .Z(n11531) );
  OR2 U7856 ( .A(n11532), .B(reset_to_pma_tx), .Z(U160_Z_0) );
  AN2 U7857 ( .A(n3179), .B(U160_DATA2_0), .Z(n11532) );
  IV U7858 ( .A(n4921), .Z(U160_DATA2_3) );
  OR2 U7859 ( .A(n3248), .B(n11533), .Z(n4921) );
  AN2 U7860 ( .A(n11534), .B(n11535), .Z(n11533) );
  OR2 U7861 ( .A(n11536), .B(n11537), .Z(n11535) );
  IV U7862 ( .A(tx_fifo_pop_pre), .Z(n11537) );
  AN2 U7863 ( .A(n11538), .B(n11539), .Z(n11536) );
  OR2 U7864 ( .A(n3250), .B(n11540), .Z(n11539) );
  AN2 U7865 ( .A(n11541), .B(n11542), .Z(n11540) );
  IV U7866 ( .A(n3252), .Z(n11541) );
  IV U7867 ( .A(n3476), .Z(n11534) );
  OR2 U7868 ( .A(n11543), .B(n11544), .Z(U160_DATA2_2) );
  OR2 U7869 ( .A(n11545), .B(n11546), .Z(n11544) );
  AN2 U7870 ( .A(n11547), .B(n3252), .Z(n11545) );
  AN2 U7871 ( .A(n11548), .B(n11542), .Z(n11547) );
  IV U7872 ( .A(n3251), .Z(n11542) );
  OR2 U7873 ( .A(n11549), .B(n11550), .Z(U160_DATA2_1) );
  OR2 U7874 ( .A(n11551), .B(n11546), .Z(n11550) );
  OR2 U7875 ( .A(n11552), .B(n3248), .Z(n11546) );
  AN2 U7876 ( .A(n3250), .B(n11548), .Z(n11552) );
  AN2 U7877 ( .A(n3251), .B(n11548), .Z(n11551) );
  OR2 U7878 ( .A(n3476), .B(n11553), .Z(n11549) );
  OR2 U7879 ( .A(n11554), .B(n11553), .Z(U160_DATA2_0) );
  AN2 U7880 ( .A(n11555), .B(n11556), .Z(n11553) );
  AN2 U7881 ( .A(n11548), .B(n3253), .Z(n11556) );
  AN2 U7882 ( .A(n11538), .B(tx_fifo_pop_pre), .Z(n11548) );
  IV U7883 ( .A(n3249), .Z(n11538) );
  AN2 U7884 ( .A(n11557), .B(n11558), .Z(n11555) );
  IV U7885 ( .A(n11559), .Z(n11558) );
  AN2 U7886 ( .A(n11560), .B(n11557), .Z(n11554) );
  IV U7887 ( .A(n3248), .Z(n11557) );
  OR2 U7888 ( .A(n11561), .B(n11543), .Z(n11560) );
  OR2 U7889 ( .A(n11562), .B(n3476), .Z(n11543) );
  IV U7890 ( .A(n11563), .Z(n11562) );
  OR2 U7891 ( .A(n11564), .B(n11559), .Z(n11563) );
  OR2 U7892 ( .A(n3250), .B(n11565), .Z(n11559) );
  OR2 U7893 ( .A(n3252), .B(n3251), .Z(n11565) );
  OR2 U7894 ( .A(n3249), .B(n3253), .Z(n11564) );
  AN2 U7895 ( .A(n3249), .B(tx_fifo_pop_pre), .Z(n11561) );
  AN2 U7896 ( .A(n10092), .B(U162_DATA3_48), .Z(U159_Z_7) );
  AN2 U7897 ( .A(n10092), .B(U162_DATA3_40), .Z(U159_Z_6) );
  OR2 U7898 ( .A(U162_DATA3_34), .B(n11566), .Z(U159_Z_5) );
  AN2 U7899 ( .A(n10092), .B(U162_DATA3_32), .Z(U159_Z_4) );
  AN2 U7900 ( .A(n10092), .B(U162_DATA3_16), .Z(U159_Z_3) );
  AN2 U7901 ( .A(n10092), .B(U162_DATA3_8), .Z(U159_Z_2) );
  OR2 U7902 ( .A(U162_DATA3_2), .B(n11566), .Z(U159_Z_1) );
  OR2 U7903 ( .A(n11567), .B(n11568), .Z(n11566) );
  OR2 U7904 ( .A(n5458), .B(n5457), .Z(n11568) );
  AN2 U7905 ( .A(n10092), .B(U162_DATA3_0), .Z(U159_Z_0) );
  OR2 U7906 ( .A(n11569), .B(n4170), .Z(U158_Z_9) );
  AN2 U7907 ( .A(U162_DATA3_41), .B(n10092), .Z(n11569) );
  OR2 U7908 ( .A(n11570), .B(n4170), .Z(U158_Z_8) );
  AN2 U7909 ( .A(U162_DATA3_33), .B(n10092), .Z(n11570) );
  OR2 U7910 ( .A(n11571), .B(n4170), .Z(U158_Z_6) );
  AN2 U7911 ( .A(U162_DATA3_25), .B(n10092), .Z(n11571) );
  OR2 U7912 ( .A(n5458), .B(n11572), .Z(U158_Z_5) );
  AN2 U7913 ( .A(U162_DATA3_24), .B(n10092), .Z(n11572) );
  OR2 U7914 ( .A(n11573), .B(n4170), .Z(U158_Z_3) );
  AN2 U7915 ( .A(U162_DATA3_17), .B(n10092), .Z(n11573) );
  OR2 U7916 ( .A(n11574), .B(n4170), .Z(U158_Z_14) );
  AN2 U7917 ( .A(U162_DATA3_57), .B(n10092), .Z(n11574) );
  OR2 U7918 ( .A(n5458), .B(n11575), .Z(U158_Z_13) );
  AN2 U7919 ( .A(U162_DATA3_56), .B(n10092), .Z(n11575) );
  IV U7920 ( .A(n3286), .Z(n5458) );
  OR2 U7921 ( .A(n11576), .B(n4170), .Z(U158_Z_11) );
  AN2 U7922 ( .A(U162_DATA3_49), .B(n10092), .Z(n11576) );
  OR2 U7923 ( .A(n11577), .B(n4170), .Z(U158_Z_1) );
  AN2 U7924 ( .A(U162_DATA3_9), .B(n10092), .Z(n11577) );
  OR2 U7925 ( .A(n11578), .B(n4170), .Z(U158_Z_0) );
  AN2 U7926 ( .A(U162_DATA3_1), .B(n10092), .Z(n11578) );
  OR2 U7927 ( .A(n11579), .B(n4172), .Z(U157_Z_5) );
  AN2 U7928 ( .A(U162_DATA3_39), .B(n10092), .Z(n11579) );
  OR2 U7929 ( .A(n11580), .B(n4172), .Z(U157_Z_4) );
  AN2 U7930 ( .A(U162_DATA3_36), .B(n10092), .Z(n11580) );
  OR2 U7931 ( .A(n11581), .B(n4172), .Z(U157_Z_3) );
  AN2 U7932 ( .A(U162_DATA3_35), .B(n10092), .Z(n11581) );
  OR2 U7933 ( .A(n11582), .B(n4172), .Z(U157_Z_2) );
  AN2 U7934 ( .A(U162_DATA3_7), .B(n10092), .Z(n11582) );
  OR2 U7935 ( .A(n11583), .B(n4172), .Z(U157_Z_1) );
  AN2 U7936 ( .A(U162_DATA3_4), .B(n10092), .Z(n11583) );
  OR2 U7937 ( .A(n11584), .B(n4172), .Z(U157_Z_0) );
  AN2 U7938 ( .A(U162_DATA3_3), .B(n10092), .Z(n11584) );
  AN2 U7939 ( .A(n11585), .B(n3284), .Z(U157_CONTROL2) );
  AN2 U7940 ( .A(n3286), .B(n11567), .Z(n11585) );
  IV U7941 ( .A(n3279), .Z(n11567) );
  OR2 U7942 ( .A(n11586), .B(n5457), .Z(U156_Z_9) );
  AN2 U7943 ( .A(U162_DATA3_21), .B(n10092), .Z(n11586) );
  OR2 U7944 ( .A(n11587), .B(n5457), .Z(U156_Z_8) );
  AN2 U7945 ( .A(U162_DATA3_20), .B(n10092), .Z(n11587) );
  OR2 U7946 ( .A(n11588), .B(n5457), .Z(U156_Z_7) );
  AN2 U7947 ( .A(U162_DATA3_19), .B(n10092), .Z(n11588) );
  OR2 U7948 ( .A(n11589), .B(n5457), .Z(U156_Z_6) );
  AN2 U7949 ( .A(U162_DATA3_15), .B(n10092), .Z(n11589) );
  OR2 U7950 ( .A(n11590), .B(n5457), .Z(U156_Z_5) );
  AN2 U7951 ( .A(U162_DATA3_14), .B(n10092), .Z(n11590) );
  OR2 U7952 ( .A(n11591), .B(n5457), .Z(U156_Z_4) );
  AN2 U7953 ( .A(U162_DATA3_13), .B(n10092), .Z(n11591) );
  OR2 U7954 ( .A(n11592), .B(n5457), .Z(U156_Z_33) );
  AN2 U7955 ( .A(U162_DATA3_63), .B(n10092), .Z(n11592) );
  OR2 U7956 ( .A(n11593), .B(n5457), .Z(U156_Z_32) );
  AN2 U7957 ( .A(U162_DATA3_62), .B(n10092), .Z(n11593) );
  OR2 U7958 ( .A(n11594), .B(n5457), .Z(U156_Z_31) );
  AN2 U7959 ( .A(U162_DATA3_61), .B(n10092), .Z(n11594) );
  OR2 U7960 ( .A(n11595), .B(n5457), .Z(U156_Z_30) );
  AN2 U7961 ( .A(U162_DATA3_60), .B(n10092), .Z(n11595) );
  OR2 U7962 ( .A(n11596), .B(n5457), .Z(U156_Z_3) );
  AN2 U7963 ( .A(U162_DATA3_12), .B(n10092), .Z(n11596) );
  OR2 U7964 ( .A(n11597), .B(n5457), .Z(U156_Z_29) );
  AN2 U7965 ( .A(U162_DATA3_59), .B(n10092), .Z(n11597) );
  OR2 U7966 ( .A(n11598), .B(n5457), .Z(U156_Z_28) );
  AN2 U7967 ( .A(U162_DATA3_55), .B(n10092), .Z(n11598) );
  OR2 U7968 ( .A(n11599), .B(n5457), .Z(U156_Z_27) );
  AN2 U7969 ( .A(U162_DATA3_54), .B(n10092), .Z(n11599) );
  OR2 U7970 ( .A(n11600), .B(n5457), .Z(U156_Z_26) );
  AN2 U7971 ( .A(U162_DATA3_53), .B(n10092), .Z(n11600) );
  OR2 U7972 ( .A(n11601), .B(n5457), .Z(U156_Z_25) );
  AN2 U7973 ( .A(U162_DATA3_52), .B(n10092), .Z(n11601) );
  OR2 U7974 ( .A(n11602), .B(n5457), .Z(U156_Z_24) );
  AN2 U7975 ( .A(U162_DATA3_51), .B(n10092), .Z(n11602) );
  OR2 U7976 ( .A(n11603), .B(n5457), .Z(U156_Z_23) );
  AN2 U7977 ( .A(U162_DATA3_47), .B(n10092), .Z(n11603) );
  OR2 U7978 ( .A(n11604), .B(n5457), .Z(U156_Z_22) );
  AN2 U7979 ( .A(U162_DATA3_46), .B(n10092), .Z(n11604) );
  OR2 U7980 ( .A(n11605), .B(n5457), .Z(U156_Z_21) );
  AN2 U7981 ( .A(U162_DATA3_45), .B(n10092), .Z(n11605) );
  OR2 U7982 ( .A(n11606), .B(n5457), .Z(U156_Z_20) );
  AN2 U7983 ( .A(U162_DATA3_44), .B(n10092), .Z(n11606) );
  OR2 U7984 ( .A(n11607), .B(n5457), .Z(U156_Z_2) );
  AN2 U7985 ( .A(U162_DATA3_11), .B(n10092), .Z(n11607) );
  OR2 U7986 ( .A(n11608), .B(n5457), .Z(U156_Z_19) );
  AN2 U7987 ( .A(U162_DATA3_43), .B(n10092), .Z(n11608) );
  OR2 U7988 ( .A(n11609), .B(n5457), .Z(U156_Z_18) );
  AN2 U7989 ( .A(U162_DATA3_38), .B(n10092), .Z(n11609) );
  OR2 U7990 ( .A(n11610), .B(n5457), .Z(U156_Z_17) );
  AN2 U7991 ( .A(U162_DATA3_37), .B(n10092), .Z(n11610) );
  OR2 U7992 ( .A(n11611), .B(n5457), .Z(U156_Z_16) );
  AN2 U7993 ( .A(U162_DATA3_31), .B(n10092), .Z(n11611) );
  OR2 U7994 ( .A(n11612), .B(n5457), .Z(U156_Z_15) );
  AN2 U7995 ( .A(U162_DATA3_30), .B(n10092), .Z(n11612) );
  OR2 U7996 ( .A(n11613), .B(n5457), .Z(U156_Z_14) );
  AN2 U7997 ( .A(U162_DATA3_29), .B(n10092), .Z(n11613) );
  OR2 U7998 ( .A(n11614), .B(n5457), .Z(U156_Z_13) );
  AN2 U7999 ( .A(U162_DATA3_28), .B(n10092), .Z(n11614) );
  OR2 U8000 ( .A(n11615), .B(n5457), .Z(U156_Z_12) );
  AN2 U8001 ( .A(U162_DATA3_27), .B(n10092), .Z(n11615) );
  OR2 U8002 ( .A(n11616), .B(n5457), .Z(U156_Z_11) );
  AN2 U8003 ( .A(U162_DATA3_23), .B(n10092), .Z(n11616) );
  OR2 U8004 ( .A(n11617), .B(n5457), .Z(U156_Z_10) );
  AN2 U8005 ( .A(U162_DATA3_22), .B(n10092), .Z(n11617) );
  OR2 U8006 ( .A(n11618), .B(n5457), .Z(U156_Z_1) );
  AN2 U8007 ( .A(U162_DATA3_6), .B(n10092), .Z(n11618) );
  OR2 U8008 ( .A(n11619), .B(n5457), .Z(U156_Z_0) );
  AN2 U8009 ( .A(n8701), .B(n3286), .Z(n5457) );
  AN2 U8010 ( .A(U162_DATA3_5), .B(n10092), .Z(n11619) );
  AN2 U8011 ( .A(n3284), .B(n11620), .Z(n10092) );
  AN2 U8012 ( .A(n3286), .B(n3279), .Z(n11620) );
  OR2 U8013 ( .A(U161_DATA3_4), .B(n11621), .Z(U155_Z_1) );
  OR2 U8014 ( .A(U161_DATA3_0), .B(n11621), .Z(U155_Z_0) );
  IV U8015 ( .A(n11622), .Z(n11621) );
  OR2 U8016 ( .A(n11623), .B(n4173), .Z(U154_Z_5) );
  AN2 U8017 ( .A(U161_DATA3_7), .B(n11622), .Z(n11623) );
  OR2 U8018 ( .A(n11624), .B(n4173), .Z(U154_Z_4) );
  AN2 U8019 ( .A(U161_DATA3_6), .B(n11622), .Z(n11624) );
  OR2 U8020 ( .A(n11625), .B(n4173), .Z(U154_Z_3) );
  AN2 U8021 ( .A(U161_DATA3_5), .B(n11622), .Z(n11625) );
  OR2 U8022 ( .A(n11626), .B(n4173), .Z(U154_Z_2) );
  AN2 U8023 ( .A(U161_DATA3_3), .B(n11622), .Z(n11626) );
  OR2 U8024 ( .A(n11627), .B(n4173), .Z(U154_Z_1) );
  AN2 U8025 ( .A(U161_DATA3_2), .B(n11622), .Z(n11627) );
  OR2 U8026 ( .A(n11628), .B(n4173), .Z(U154_Z_0) );
  AN2 U8027 ( .A(U161_DATA3_1), .B(n11622), .Z(n11628) );
  AN2 U8028 ( .A(n3290), .B(n11629), .Z(n11622) );
  AN2 U8029 ( .A(n3281), .B(n3288), .Z(n11629) );
  AN2 U8030 ( .A(n2937), .B(n11630), .Z(U119_Z_3) );
  OR2 U8031 ( .A(n11631), .B(n11632), .Z(n11630) );
  OR2 U8032 ( .A(n11633), .B(n11634), .Z(n11632) );
  AN2 U8033 ( .A(U124_CONTROL2), .B(n11635), .Z(n11634) );
  AN2 U8034 ( .A(n4915), .B(n2953), .Z(U124_CONTROL2) );
  AN2 U8035 ( .A(U141_CONTROL2), .B(n11636), .Z(n11633) );
  AN2 U8036 ( .A(n4909), .B(n11637), .Z(U141_CONTROL2) );
  OR2 U8037 ( .A(n11638), .B(n11639), .Z(n11631) );
  OR2 U8038 ( .A(n11640), .B(n11641), .Z(n11639) );
  AN2 U8039 ( .A(n11642), .B(U150_DATA3_0), .Z(n11641) );
  AN2 U8040 ( .A(n11643), .B(n4915), .Z(n11640) );
  OR2 U8041 ( .A(n11644), .B(n11645), .Z(n11643) );
  AN2 U8042 ( .A(n11646), .B(n11647), .Z(n11644) );
  AN2 U8043 ( .A(n2974), .B(n11648), .Z(n11638) );
  AN2 U8044 ( .A(n2937), .B(n11649), .Z(U119_Z_2) );
  OR2 U8045 ( .A(n11650), .B(n11651), .Z(n11649) );
  OR2 U8046 ( .A(n11652), .B(n11653), .Z(n11651) );
  OR2 U8047 ( .A(n11654), .B(n11655), .Z(n11653) );
  AN2 U8048 ( .A(n2977), .B(n11645), .Z(n11655) );
  AN2 U8049 ( .A(n2975), .B(n11635), .Z(n11654) );
  OR2 U8050 ( .A(n11656), .B(n11657), .Z(n11650) );
  OR2 U8051 ( .A(n11658), .B(n11659), .Z(n11657) );
  AN2 U8052 ( .A(n11642), .B(U151_DATA3_0), .Z(n11659) );
  AN2 U8053 ( .A(n11648), .B(n11660), .Z(n11658) );
  OR2 U8054 ( .A(n4912), .B(n4909), .Z(n11660) );
  IV U8055 ( .A(n2968), .Z(n4909) );
  AN2 U8056 ( .A(n2979), .B(n11636), .Z(n11656) );
  AN2 U8057 ( .A(n2937), .B(n11661), .Z(U119_Z_1) );
  OR2 U8058 ( .A(n11662), .B(n11663), .Z(n11661) );
  OR2 U8059 ( .A(n11664), .B(n11665), .Z(n11663) );
  OR2 U8060 ( .A(n11666), .B(n11667), .Z(n11665) );
  AN2 U8061 ( .A(n11635), .B(n4912), .Z(n11667) );
  IV U8062 ( .A(n2953), .Z(n4912) );
  AN2 U8063 ( .A(U140_CONTROL2), .B(n11636), .Z(n11666) );
  AN2 U8064 ( .A(n2968), .B(n11668), .Z(U140_CONTROL2) );
  AN2 U8065 ( .A(n4914), .B(n11637), .Z(n11668) );
  AN2 U8066 ( .A(n2985), .B(n11645), .Z(n11664) );
  OR2 U8067 ( .A(n11669), .B(n11670), .Z(n11662) );
  OR2 U8068 ( .A(n11671), .B(n11672), .Z(n11670) );
  AN2 U8069 ( .A(n11642), .B(U152_DATA3_0), .Z(n11672) );
  AN2 U8070 ( .A(n11673), .B(n4916), .Z(n11671) );
  AN2 U8071 ( .A(n2987), .B(n11648), .Z(n11669) );
  AN2 U8072 ( .A(n2937), .B(n11674), .Z(U119_Z_0) );
  OR2 U8073 ( .A(n11675), .B(n11676), .Z(n11674) );
  OR2 U8074 ( .A(n11677), .B(n11678), .Z(n11676) );
  OR2 U8075 ( .A(n11679), .B(n11680), .Z(n11677) );
  AN2 U8076 ( .A(n2988), .B(n11635), .Z(n11680) );
  AN2 U8077 ( .A(n2972), .B(n11636), .Z(n11679) );
  OR2 U8078 ( .A(n11681), .B(n11682), .Z(n11675) );
  OR2 U8079 ( .A(n11683), .B(n11684), .Z(n11682) );
  AN2 U8080 ( .A(n11648), .B(n4914), .Z(n11684) );
  IV U8081 ( .A(n2958), .Z(n4914) );
  AN2 U8082 ( .A(n11642), .B(U153_DATA2_0), .Z(n11683) );
  OR2 U8083 ( .A(n11685), .B(n11686), .Z(n11681) );
  AN2 U8084 ( .A(n11687), .B(n4916), .Z(n11686) );
  AN2 U8085 ( .A(n11688), .B(n4915), .Z(n11685) );
  IV U8086 ( .A(n2961), .Z(n4915) );
  OR2 U8087 ( .A(n11648), .B(n11687), .Z(n11688) );
  AN2 U8088 ( .A(n2937), .B(n11689), .Z(U118_Z_1) );
  OR2 U8089 ( .A(n11690), .B(n11678), .Z(n11689) );
  OR2 U8090 ( .A(n11691), .B(n11652), .Z(n11678) );
  OR2 U8091 ( .A(n11692), .B(n11693), .Z(n11652) );
  AN2 U8092 ( .A(n2884), .B(n11646), .Z(n11693) );
  AN2 U8093 ( .A(n2915), .B(n11648), .Z(n11692) );
  AN2 U8094 ( .A(n2892), .B(n11645), .Z(n11691) );
  OR2 U8095 ( .A(n11694), .B(n11695), .Z(n11690) );
  OR2 U8096 ( .A(n11696), .B(n11697), .Z(n11695) );
  AN2 U8097 ( .A(n2900), .B(n11636), .Z(n11697) );
  AN2 U8098 ( .A(n11642), .B(U148_DATA3_0), .Z(n11696) );
  AN2 U8099 ( .A(U122_CONTROL2), .B(n11635), .Z(n11694) );
  AN2 U8100 ( .A(n2923), .B(n11698), .Z(U122_CONTROL2) );
  OR2 U8101 ( .A(n11699), .B(reset_to_pma_tx), .Z(U118_Z_0) );
  AN2 U8102 ( .A(n11700), .B(n2937), .Z(n11699) );
  AN2 U8103 ( .A(n11642), .B(U149_DATA2_0), .Z(n11700) );
  OR2 U8104 ( .A(n11701), .B(n11702), .Z(n11642) );
  OR2 U8105 ( .A(n11703), .B(n11704), .Z(n11702) );
  AN2 U8106 ( .A(n11673), .B(n2948), .Z(n11704) );
  AN2 U8107 ( .A(n11646), .B(n11705), .Z(n11673) );
  AN2 U8108 ( .A(n11647), .B(n2961), .Z(n11705) );
  IV U8109 ( .A(n2884), .Z(n11647) );
  AN2 U8110 ( .A(n11698), .B(n11706), .Z(n11703) );
  OR2 U8111 ( .A(n11707), .B(n11708), .Z(n11706) );
  OR2 U8112 ( .A(n11709), .B(n11710), .Z(n11708) );
  AN2 U8113 ( .A(n11711), .B(n11645), .Z(n11710) );
  IV U8114 ( .A(n11712), .Z(n11711) );
  OR2 U8115 ( .A(n4916), .B(n2892), .Z(n11712) );
  IV U8116 ( .A(n2948), .Z(n4916) );
  AN2 U8117 ( .A(n11713), .B(n11714), .Z(n11709) );
  AN2 U8118 ( .A(n2958), .B(n11715), .Z(n11714) );
  IV U8119 ( .A(n2915), .Z(n11715) );
  AN2 U8120 ( .A(n11648), .B(n2968), .Z(n11713) );
  IV U8121 ( .A(n11716), .Z(n11648) );
  AN2 U8122 ( .A(n11635), .B(n11717), .Z(n11707) );
  IV U8123 ( .A(n2923), .Z(n11717) );
  IV U8124 ( .A(n11718), .Z(n11635) );
  AN2 U8125 ( .A(n2953), .B(n2961), .Z(n11698) );
  OR2 U8126 ( .A(n11719), .B(n11720), .Z(n11701) );
  AN2 U8127 ( .A(n11721), .B(n11636), .Z(n11720) );
  IV U8128 ( .A(n11722), .Z(n11636) );
  AN2 U8129 ( .A(n11723), .B(n2968), .Z(n11721) );
  AN2 U8130 ( .A(n2958), .B(n11637), .Z(n11723) );
  IV U8131 ( .A(n2900), .Z(n11637) );
  AN2 U8132 ( .A(n11724), .B(n11722), .Z(n11719) );
  OR2 U8133 ( .A(n2867), .B(n2868), .Z(n11722) );
  AN2 U8134 ( .A(n11725), .B(n11726), .Z(n11724) );
  IV U8135 ( .A(n11687), .Z(n11726) );
  OR2 U8136 ( .A(n11646), .B(n11645), .Z(n11687) );
  IV U8137 ( .A(n11727), .Z(n11645) );
  AN2 U8138 ( .A(n11728), .B(n11729), .Z(n11727) );
  OR2 U8139 ( .A(n2863), .B(n2864), .Z(n11729) );
  OR2 U8140 ( .A(n2871), .B(n2872), .Z(n11728) );
  AN2 U8141 ( .A(n2862), .B(n2861), .Z(n11646) );
  AN2 U8142 ( .A(n11716), .B(n11718), .Z(n11725) );
  OR2 U8143 ( .A(n2879), .B(n2880), .Z(n11718) );
  OR2 U8144 ( .A(n2875), .B(n2876), .Z(n11716) );
  OR2 U8145 ( .A(n11730), .B(n11731), .Z(U117_Z_9) );
  AN2 U8146 ( .A(n11732), .B(n11733), .Z(n11731) );
  AN2 U8147 ( .A(n11734), .B(n11735), .Z(n11732) );
  AN2 U8148 ( .A(U3_U1_DATA1_9), .B(n11736), .Z(n11730) );
  OR2 U8149 ( .A(n11737), .B(n11738), .Z(U117_Z_8) );
  AN2 U8150 ( .A(n11739), .B(n11740), .Z(n11738) );
  AN2 U8151 ( .A(n11741), .B(n11734), .Z(n11739) );
  AN2 U8152 ( .A(n11742), .B(U3_U1_DATA1_7), .Z(n11741) );
  AN2 U8153 ( .A(U3_U1_DATA1_8), .B(n11743), .Z(n11737) );
  OR2 U8154 ( .A(n11744), .B(n11745), .Z(n11743) );
  AN2 U8155 ( .A(n11746), .B(n11747), .Z(n11744) );
  OR2 U8156 ( .A(n11748), .B(n11749), .Z(U117_Z_7) );
  AN2 U8157 ( .A(n11750), .B(n11747), .Z(n11749) );
  AN2 U8158 ( .A(n11734), .B(n11742), .Z(n11750) );
  IV U8159 ( .A(n11751), .Z(n11742) );
  AN2 U8160 ( .A(U3_U1_DATA1_7), .B(n11745), .Z(n11748) );
  OR2 U8161 ( .A(n11752), .B(n11753), .Z(n11745) );
  AN2 U8162 ( .A(n11746), .B(n11751), .Z(n11752) );
  OR2 U8163 ( .A(n11754), .B(n11755), .Z(U117_Z_6) );
  AN2 U8164 ( .A(n11756), .B(n11757), .Z(n11755) );
  AN2 U8165 ( .A(n11758), .B(n11734), .Z(n11756) );
  AN2 U8166 ( .A(n11759), .B(U3_U1_DATA1_5), .Z(n11758) );
  AN2 U8167 ( .A(U3_U1_DATA1_6), .B(n11760), .Z(n11754) );
  OR2 U8168 ( .A(n11761), .B(n11762), .Z(n11760) );
  AN2 U8169 ( .A(n11746), .B(n11763), .Z(n11761) );
  OR2 U8170 ( .A(n11764), .B(n11765), .Z(U117_Z_5) );
  AN2 U8171 ( .A(n11766), .B(n11763), .Z(n11765) );
  AN2 U8172 ( .A(n11734), .B(n11759), .Z(n11766) );
  IV U8173 ( .A(n11767), .Z(n11759) );
  AN2 U8174 ( .A(U3_U1_DATA1_5), .B(n11762), .Z(n11764) );
  OR2 U8175 ( .A(n11768), .B(n11753), .Z(n11762) );
  AN2 U8176 ( .A(n11746), .B(n11767), .Z(n11768) );
  OR2 U8177 ( .A(n11769), .B(n11770), .Z(U117_Z_4) );
  AN2 U8178 ( .A(n11771), .B(n11772), .Z(n11770) );
  AN2 U8179 ( .A(n11773), .B(n11734), .Z(n11771) );
  AN2 U8180 ( .A(n11774), .B(U3_U1_DATA1_3), .Z(n11773) );
  AN2 U8181 ( .A(U3_U1_DATA1_4), .B(n11775), .Z(n11769) );
  OR2 U8182 ( .A(n11776), .B(n11777), .Z(n11775) );
  AN2 U8183 ( .A(n11746), .B(n11778), .Z(n11776) );
  OR2 U8184 ( .A(n11779), .B(n11780), .Z(U117_Z_3) );
  AN2 U8185 ( .A(n11781), .B(n11778), .Z(n11780) );
  AN2 U8186 ( .A(n11734), .B(n11774), .Z(n11781) );
  IV U8187 ( .A(n11782), .Z(n11774) );
  AN2 U8188 ( .A(U3_U1_DATA1_3), .B(n11777), .Z(n11779) );
  OR2 U8189 ( .A(n11783), .B(n11753), .Z(n11777) );
  AN2 U8190 ( .A(n11746), .B(n11782), .Z(n11783) );
  OR2 U8191 ( .A(n11784), .B(n11785), .Z(U117_Z_2) );
  AN2 U8192 ( .A(n11786), .B(n11787), .Z(n11785) );
  AN2 U8193 ( .A(n11788), .B(n11734), .Z(n11786) );
  AN2 U8194 ( .A(U3_U1_DATA1_1), .B(U3_U1_DATA1_0), .Z(n11788) );
  AN2 U8195 ( .A(U3_U1_DATA1_2), .B(n11789), .Z(n11784) );
  OR2 U8196 ( .A(n11790), .B(n11791), .Z(n11789) );
  AN2 U8197 ( .A(n11746), .B(n11792), .Z(n11790) );
  OR2 U8198 ( .A(n11793), .B(n11794), .Z(U117_Z_15) );
  AN2 U8199 ( .A(n11795), .B(n11796), .Z(n11794) );
  IV U8200 ( .A(U3_U1_DATA1_15), .Z(n11796) );
  AN2 U8201 ( .A(n11797), .B(U3_U1_DATA1_14), .Z(n11795) );
  AN2 U8202 ( .A(U3_U1_DATA1_15), .B(n11798), .Z(n11793) );
  OR2 U8203 ( .A(n11799), .B(n11800), .Z(n11798) );
  AN2 U8204 ( .A(n11746), .B(n11801), .Z(n11799) );
  OR2 U8205 ( .A(n11802), .B(n11803), .Z(U117_Z_14) );
  AN2 U8206 ( .A(U3_U1_DATA1_14), .B(n11800), .Z(n11803) );
  OR2 U8207 ( .A(n11804), .B(n11805), .Z(n11800) );
  AN2 U8208 ( .A(n11746), .B(n11806), .Z(n11804) );
  AN2 U8209 ( .A(n11797), .B(n11801), .Z(n11802) );
  IV U8210 ( .A(U3_U1_DATA1_14), .Z(n11801) );
  AN2 U8211 ( .A(n11807), .B(n11808), .Z(n11797) );
  AN2 U8212 ( .A(U3_U1_DATA1_13), .B(n11734), .Z(n11808) );
  OR2 U8213 ( .A(n11809), .B(n11810), .Z(U117_Z_13) );
  AN2 U8214 ( .A(n11811), .B(n11806), .Z(n11810) );
  IV U8215 ( .A(U3_U1_DATA1_13), .Z(n11806) );
  AN2 U8216 ( .A(n11807), .B(n11734), .Z(n11811) );
  IV U8217 ( .A(n11812), .Z(n11807) );
  AN2 U8218 ( .A(U3_U1_DATA1_13), .B(n11805), .Z(n11809) );
  OR2 U8219 ( .A(n11813), .B(n11753), .Z(n11805) );
  AN2 U8220 ( .A(n11746), .B(n11812), .Z(n11813) );
  OR2 U8221 ( .A(n11814), .B(n11815), .Z(n11812) );
  OR2 U8222 ( .A(n11816), .B(n11817), .Z(n11815) );
  OR2 U8223 ( .A(n11818), .B(n11819), .Z(U117_Z_12) );
  AN2 U8224 ( .A(n11820), .B(n11816), .Z(n11819) );
  IV U8225 ( .A(U3_U1_DATA1_12), .Z(n11816) );
  AN2 U8226 ( .A(n11821), .B(n11822), .Z(n11820) );
  AN2 U8227 ( .A(n11734), .B(U3_U1_DATA1_11), .Z(n11821) );
  AN2 U8228 ( .A(U3_U1_DATA1_12), .B(n11823), .Z(n11818) );
  OR2 U8229 ( .A(n11824), .B(n11825), .Z(n11823) );
  AN2 U8230 ( .A(n11746), .B(n11817), .Z(n11824) );
  OR2 U8231 ( .A(n11826), .B(n11827), .Z(U117_Z_11) );
  AN2 U8232 ( .A(n11828), .B(n11817), .Z(n11827) );
  IV U8233 ( .A(U3_U1_DATA1_11), .Z(n11817) );
  AN2 U8234 ( .A(n11822), .B(n11734), .Z(n11828) );
  IV U8235 ( .A(n11814), .Z(n11822) );
  AN2 U8236 ( .A(U3_U1_DATA1_11), .B(n11825), .Z(n11826) );
  OR2 U8237 ( .A(n11829), .B(n11753), .Z(n11825) );
  AN2 U8238 ( .A(n11746), .B(n11814), .Z(n11829) );
  OR2 U8239 ( .A(n11830), .B(n11831), .Z(n11814) );
  OR2 U8240 ( .A(n11733), .B(n11832), .Z(n11831) );
  OR2 U8241 ( .A(n11833), .B(n11834), .Z(U117_Z_10) );
  AN2 U8242 ( .A(n11835), .B(n11832), .Z(n11834) );
  IV U8243 ( .A(U3_U1_DATA1_10), .Z(n11832) );
  AN2 U8244 ( .A(n11836), .B(n11734), .Z(n11835) );
  AN2 U8245 ( .A(n11735), .B(U3_U1_DATA1_9), .Z(n11836) );
  IV U8246 ( .A(n11830), .Z(n11735) );
  AN2 U8247 ( .A(U3_U1_DATA1_10), .B(n11837), .Z(n11833) );
  OR2 U8248 ( .A(n11838), .B(n11736), .Z(n11837) );
  OR2 U8249 ( .A(n11839), .B(n11753), .Z(n11736) );
  AN2 U8250 ( .A(n11746), .B(n11830), .Z(n11839) );
  OR2 U8251 ( .A(n11751), .B(n11840), .Z(n11830) );
  OR2 U8252 ( .A(n11740), .B(n11747), .Z(n11840) );
  IV U8253 ( .A(U3_U1_DATA1_7), .Z(n11747) );
  IV U8254 ( .A(U3_U1_DATA1_8), .Z(n11740) );
  OR2 U8255 ( .A(n11767), .B(n11841), .Z(n11751) );
  OR2 U8256 ( .A(n11757), .B(n11763), .Z(n11841) );
  IV U8257 ( .A(U3_U1_DATA1_5), .Z(n11763) );
  IV U8258 ( .A(U3_U1_DATA1_6), .Z(n11757) );
  OR2 U8259 ( .A(n11782), .B(n11842), .Z(n11767) );
  OR2 U8260 ( .A(n11772), .B(n11778), .Z(n11842) );
  IV U8261 ( .A(U3_U1_DATA1_3), .Z(n11778) );
  IV U8262 ( .A(U3_U1_DATA1_4), .Z(n11772) );
  OR2 U8263 ( .A(n11792), .B(n11843), .Z(n11782) );
  OR2 U8264 ( .A(n11844), .B(n11787), .Z(n11843) );
  IV U8265 ( .A(U3_U1_DATA1_2), .Z(n11787) );
  AN2 U8266 ( .A(n11746), .B(n11733), .Z(n11838) );
  IV U8267 ( .A(U3_U1_DATA1_9), .Z(n11733) );
  OR2 U8268 ( .A(n11845), .B(n11846), .Z(U117_Z_1) );
  AN2 U8269 ( .A(n11847), .B(n11792), .Z(n11846) );
  IV U8270 ( .A(U3_U1_DATA1_1), .Z(n11792) );
  AN2 U8271 ( .A(n11734), .B(U3_U1_DATA1_0), .Z(n11847) );
  AN2 U8272 ( .A(U3_U1_DATA1_1), .B(n11791), .Z(n11845) );
  OR2 U8273 ( .A(n11848), .B(n11753), .Z(n11791) );
  AN2 U8274 ( .A(n11746), .B(n11844), .Z(n11848) );
  OR2 U8275 ( .A(n11849), .B(n11850), .Z(U117_Z_0) );
  AN2 U8276 ( .A(n11753), .B(U3_U1_DATA1_0), .Z(n11850) );
  AN2 U8277 ( .A(n11746), .B(n2689), .Z(n11753) );
  IV U8278 ( .A(n11851), .Z(n11746) );
  AN2 U8279 ( .A(n11734), .B(n11844), .Z(n11849) );
  IV U8280 ( .A(U3_U1_DATA1_0), .Z(n11844) );
  IV U8281 ( .A(n11852), .Z(n11734) );
  OR2 U8282 ( .A(n2689), .B(n11851), .Z(n11852) );
  OR2 U8283 ( .A(n8999), .B(n9011), .Z(n11851) );
  AN2 U8284 ( .A(n9050), .B(U72_DATA3_0), .Z(n9011) );
  IV U8285 ( .A(n11853), .Z(n9050) );
  OR2 U8286 ( .A(n2541), .B(n2540), .Z(n11853) );
  AN2 U8287 ( .A(U71_DATA3_0), .B(n8719), .Z(n8999) );
  IV U8288 ( .A(n9043), .Z(n8719) );
  OR2 U8289 ( .A(n2544), .B(n2545), .Z(n9043) );
endmodule

