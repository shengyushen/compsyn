
module PCIEXP_TX ( PCLK250, RST_BeaconEnable_R0, CNTL_RESETN_P0, 
        CNTL_Loopback_P0, CNTL_TXEnable_P0, RX_LoopbackData_P2, TXCOMPLIANCE, 
        TXDATA, TXDATAK, TXELECIDLE, HSS_TXBEACONCMD, HSS_TXD, HSS_TXELECIDLE
 );
  input [9:0] RX_LoopbackData_P2;
  input [7:0] TXDATA;
  output [9:0] HSS_TXD;
  input PCLK250, RST_BeaconEnable_R0, CNTL_RESETN_P0, CNTL_Loopback_P0,
         CNTL_TXEnable_P0, TXCOMPLIANCE, TXDATAK, TXELECIDLE;
  output HSS_TXBEACONCMD, HSS_TXELECIDLE;
  wire   n3, n4, n10, n11, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n25, n26, n28, n29, n30, n31, n32, n33, n35, n36, n37, n39, n40, n41,
         n44, n46, n48, n49, n52, n55, n58, n59, n60, n63, n64, n65, n68, n69,
         n71, n72, n73, n74, n76, n78, n80, n82, n84, n86, n87, n89, n91, n93,
         n94, n96, n97, n98, n100, n101, n102, n104, n105, n106, n108, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n140, n141, n142, n145, n146, n147,
         n148, n149, n150, n151, n153, n154, n157, n158, n159, n160, n162,
         n163, n164, n165, n166, n167, n168, n181, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, U6_Z_0, U6_DATA2_0,
         U5_DATA2_4, U5_DATA2_5, U4_Z_0, n325, n327, n328, n330, n332, n334,
         n336, n338, n340, n342, n344, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540;
  wire   [5:9] n;

  OR2 C36 ( .A(n400), .B(n401), .Z(n25) );
  OR2 C37 ( .A(n204), .B(n25), .Z(n26) );
  AN2 C39 ( .A(n198), .B(n197), .Z(n28) );
  AN2 C40 ( .A(n199), .B(n28), .Z(n29) );
  AN2 C41 ( .A(n200), .B(n29), .Z(n30) );
  OR2 C42 ( .A(n198), .B(n197), .Z(n31) );
  OR2 C43 ( .A(n199), .B(n31), .Z(n32) );
  OR2 C44 ( .A(n200), .B(n32), .Z(n33) );
  AN2 C46 ( .A(n203), .B(n202), .Z(n35) );
  AN2 C47 ( .A(n204), .B(n35), .Z(n36) );
  OR2 C48 ( .A(U5_DATA2_5), .B(U5_DATA2_4), .Z(n37) );
  AN2 C50 ( .A(U5_DATA2_5), .B(U5_DATA2_4), .Z(n39) );
  OR2 C53 ( .A(n203), .B(n202), .Z(n40) );
  OR2 C54 ( .A(n204), .B(n40), .Z(n41) );
  OR2 C58 ( .A(n397), .B(n40), .Z(n44) );
  OR2 C60 ( .A(n200), .B(n199), .Z(n46) );
  OR2 C67 ( .A(n420), .B(n68), .Z(n48) );
  OR2 C68 ( .A(n201), .B(n48), .Z(n49) );
  OR2 C75 ( .A(n411), .B(n69), .Z(n52) );
  OR2 C80 ( .A(n420), .B(n32), .Z(n55) );
  OR2 C83 ( .A(n198), .B(n429), .Z(n58) );
  OR2 C84 ( .A(n199), .B(n58), .Z(n59) );
  OR2 C85 ( .A(n200), .B(n59), .Z(n60) );
  OR2 C881 ( .A(n428), .B(n197), .Z(n63) );
  OR2 C891 ( .A(n199), .B(n63), .Z(n64) );
  OR2 C901 ( .A(n200), .B(n64), .Z(n65) );
  OR2 C94 ( .A(n427), .B(n31), .Z(n68) );
  OR2 C951 ( .A(n200), .B(n68), .Z(n69) );
  OR2 C100 ( .A(n428), .B(n429), .Z(n71) );
  OR2 C101 ( .A(n427), .B(n71), .Z(n72) );
  OR2 C102 ( .A(n200), .B(n72), .Z(n73) );
  OR2 C103 ( .A(n201), .B(n73), .Z(n74) );
  OR2 C108 ( .A(n201), .B(n33), .Z(n76) );
  OR2 C114 ( .A(n201), .B(n60), .Z(n78) );
  OR2 C120 ( .A(n201), .B(n65), .Z(n80) );
  OR2 C126 ( .A(n201), .B(n69), .Z(n82) );
  OR2 C132 ( .A(n201), .B(n55), .Z(n84) );
  OR2 C140 ( .A(n420), .B(n72), .Z(n86) );
  OR2 C141 ( .A(n201), .B(n86), .Z(n87) );
  OR2 C148 ( .A(n411), .B(n55), .Z(n89) );
  OR2 C154 ( .A(n411), .B(n33), .Z(n91) );
  AN2 C159 ( .A(n201), .B(n30), .Z(n93) );
  OR2 C167 ( .A(n411), .B(n73), .Z(n94) );
  OR2 C174 ( .A(n199), .B(n71), .Z(n96) );
  OR2 C175 ( .A(n420), .B(n96), .Z(n97) );
  OR2 C176 ( .A(n411), .B(n97), .Z(n98) );
  OR2 C183 ( .A(n427), .B(n58), .Z(n100) );
  OR2 C184 ( .A(n420), .B(n100), .Z(n101) );
  OR2 C185 ( .A(n411), .B(n101), .Z(n102) );
  OR2 C192 ( .A(n427), .B(n63), .Z(n104) );
  OR2 C193 ( .A(n420), .B(n104), .Z(n105) );
  OR2 C194 ( .A(n411), .B(n105), .Z(n106) );
  OR2 C202 ( .A(n411), .B(n48), .Z(n108) );
  OR2 C206 ( .A(n111), .B(n425), .Z(n[5]) );
  AN2 C207 ( .A(n198), .B(n426), .Z(n111) );
  OR2 C209 ( .A(n112), .B(n409), .Z(n[6]) );
  OR2 C210 ( .A(n199), .B(n425), .Z(n112) );
  AN2 C211 ( .A(n200), .B(n426), .Z(n[7]) );
  OR2 C213 ( .A(n113), .B(n115), .Z(n[8]) );
  OR2 C215 ( .A(n114), .B(n421), .Z(n115) );
  OR2 C216 ( .A(n423), .B(n422), .Z(n114) );
  OR2 C217 ( .A(n125), .B(n126), .Z(n[9]) );
  OR2 C218 ( .A(n124), .B(n93), .Z(n125) );
  OR2 C219 ( .A(n123), .B(n410), .Z(n124) );
  OR2 C220 ( .A(n122), .B(n419), .Z(n123) );
  OR2 C221 ( .A(n117), .B(n121), .Z(n122) );
  AN2 C222 ( .A(n424), .B(n116), .Z(n117) );
  AN2 C224 ( .A(n120), .B(n411), .Z(n121) );
  AN2 C225 ( .A(n118), .B(n119), .Z(n120) );
  AN2 C229 ( .A(n403), .B(n196), .Z(n126) );
  OR2 C230 ( .A(n131), .B(n409), .Z(n10) );
  OR2 C231 ( .A(n130), .B(n412), .Z(n131) );
  OR2 C232 ( .A(n129), .B(n413), .Z(n130) );
  OR2 C233 ( .A(n128), .B(n414), .Z(n129) );
  OR2 C234 ( .A(n127), .B(n415), .Z(n128) );
  OR2 C235 ( .A(n417), .B(n416), .Z(n127) );
  OR2 C236 ( .A(n136), .B(n137), .Z(n11) );
  OR2 C237 ( .A(n135), .B(n93), .Z(n136) );
  OR2 C238 ( .A(n134), .B(n404), .Z(n135) );
  OR2 C239 ( .A(n133), .B(n405), .Z(n134) );
  OR2 C240 ( .A(n132), .B(n406), .Z(n133) );
  OR2 C241 ( .A(n408), .B(n407), .Z(n132) );
  AN2 C242 ( .A(n403), .B(n196), .Z(n137) );
  AN2 C243 ( .A(n142), .B(n36), .Z(n13) );
  OR2 C244 ( .A(n141), .B(n196), .Z(n142) );
  OR2 C245 ( .A(n138), .B(n140), .Z(n141) );
  AN2 C246 ( .A(n393), .B(n392), .Z(n138) );
  AN2 C247 ( .A(n434), .B(n39), .Z(n140) );
  AN2 C249 ( .A(n202), .B(n391), .Z(n14) );
  OR2 C251 ( .A(n203), .B(n398), .Z(n15) );
  OR2 C252 ( .A(n145), .B(n13), .Z(n16) );
  AN2 C253 ( .A(n147), .B(n397), .Z(n145) );
  OR2 C256 ( .A(n398), .B(n396), .Z(n17) );
  AN2 C257 ( .A(n146), .B(n147), .Z(n18) );
  AN2 C258 ( .A(n403), .B(n196), .Z(n146) );
  OR2 C260 ( .A(n150), .B(n403), .Z(n19) );
  OR2 C261 ( .A(n149), .B(n404), .Z(n150) );
  OR2 C262 ( .A(n148), .B(n405), .Z(n149) );
  OR2 C263 ( .A(n407), .B(n406), .Z(n148) );
  OR2 C265 ( .A(n10), .B(n11), .Z(n151) );
  AN2 C266 ( .A(n194), .B(n154), .Z(n4) );
  OR2 C269 ( .A(n17), .B(n36), .Z(n153) );
  AN2 C270 ( .A(n395), .B(n3), .Z(n20) );
  OR2 C272 ( .A(n160), .B(n162), .Z(n21) );
  OR2 C273 ( .A(n157), .B(n159), .Z(n160) );
  AN2 C274 ( .A(n394), .B(n10), .Z(n157) );
  AN2 C276 ( .A(n20), .B(n158), .Z(n159) );
  OR2 C277 ( .A(n418), .B(n11), .Z(n158) );
  AN2 C278 ( .A(n402), .B(n196), .Z(n162) );
  OR2 C280 ( .A(n164), .B(n166), .Z(n22) );
  AN2 C281 ( .A(n434), .B(n163), .Z(n164) );
  OR2 C283 ( .A(n17), .B(n18), .Z(n163) );
  AN2 C284 ( .A(n393), .B(n165), .Z(n166) );
  OR2 C285 ( .A(n399), .B(n36), .Z(n165) );
  IV I_3 ( .A(CNTL_Loopback_P0), .Z(n181) );
  AN2 C95 ( .A(CNTL_TXEnable_P0), .B(n167), .Z(U6_DATA2_0) );
  IV I_1 ( .A(TXELECIDLE), .Z(n167) );
  AN2 C93 ( .A(RST_BeaconEnable_R0), .B(n167), .Z(HSS_TXBEACONCMD) );
  IV I_0 ( .A(CNTL_RESETN_P0), .Z(n168) );
  FD1 InputDataK_P0_reg ( .D(n390), .CP(PCLK250), .Q(n196) );
  FD1 InputCompliance_P0_reg ( .D(n389), .CP(PCLK250), .Q(n195) );
  FD1 InputData_P0_reg_7_ ( .D(n388), .CP(PCLK250), .Q(n204) );
  FD1 InputData_P0_reg_6_ ( .D(n387), .CP(PCLK250), .Q(n203) );
  FD1 InputData_P0_reg_5_ ( .D(n386), .CP(PCLK250), .Q(n202) );
  FD1 InputData_P0_reg_4_ ( .D(n385), .CP(PCLK250), .Q(n201) );
  FD1 InputData_P0_reg_3_ ( .D(n384), .CP(PCLK250), .Q(n200) );
  FD1 InputData_P0_reg_2_ ( .D(n383), .CP(PCLK250), .Q(n199) );
  FD1 InputData_P0_reg_1_ ( .D(n382), .CP(PCLK250), .Q(n198) );
  FD1 InputData_P0_reg_0_ ( .D(n381), .CP(PCLK250), .Q(n197) );
  FD1 InputDataEnable_P0_reg ( .D(U6_Z_0), .CP(PCLK250), .Q(n194) );
  FD1 OutputElecIdle_P0_reg ( .D(U4_Z_0), .CP(PCLK250), .Q(HSS_TXELECIDLE) );
  FD1 DISPARITY_P0_reg ( .D(n4), .CP(PCLK250), .Q(n3) );
  FD1 OutputData_P0_reg_7_ ( .D(n380), .CP(PCLK250), .Q(HSS_TXD[7]) );
  FD1 OutputData_P0_reg_8_ ( .D(n379), .CP(PCLK250), .Q(HSS_TXD[8]) );
  FD1 OutputData_P0_reg_4_ ( .D(n378), .CP(PCLK250), .Q(HSS_TXD[4]) );
  FD1 OutputData_P0_reg_9_ ( .D(n377), .CP(PCLK250), .Q(HSS_TXD[9]) );
  FD1 OutputData_P0_reg_6_ ( .D(n376), .CP(PCLK250), .Q(HSS_TXD[6]) );
  FD1 OutputData_P0_reg_5_ ( .D(n375), .CP(PCLK250), .Q(HSS_TXD[5]) );
  FD1 OutputData_P0_reg_0_ ( .D(n374), .CP(PCLK250), .Q(HSS_TXD[0]) );
  FD1 OutputData_P0_reg_1_ ( .D(n373), .CP(PCLK250), .Q(HSS_TXD[1]) );
  FD1 OutputData_P0_reg_2_ ( .D(n372), .CP(PCLK250), .Q(HSS_TXD[2]) );
  FD1 OutputData_P0_reg_3_ ( .D(n371), .CP(PCLK250), .Q(HSS_TXD[3]) );
  AN2 U88 ( .A(U6_DATA2_0), .B(TXDATA[0]), .Z(n325) );
  AN2 U91 ( .A(TXDATA[1]), .B(U6_DATA2_0), .Z(n328) );
  AN2 U94 ( .A(TXDATA[2]), .B(U6_DATA2_0), .Z(n330) );
  AN2 U97 ( .A(TXDATA[3]), .B(U6_DATA2_0), .Z(n332) );
  AN2 U100 ( .A(TXDATA[4]), .B(U6_DATA2_0), .Z(n334) );
  AN2 U103 ( .A(TXDATA[5]), .B(U6_DATA2_0), .Z(n336) );
  AN2 U106 ( .A(TXDATA[6]), .B(U6_DATA2_0), .Z(n338) );
  AN2 U109 ( .A(TXDATA[7]), .B(U6_DATA2_0), .Z(n340) );
  AN2 U112 ( .A(TXCOMPLIANCE), .B(U6_DATA2_0), .Z(n342) );
  IV U115 ( .A(U6_DATA2_0), .Z(n327) );
  AN2 U116 ( .A(TXDATAK), .B(U6_DATA2_0), .Z(n344) );
  AN2 U181 ( .A(CNTL_RESETN_P0), .B(U6_DATA2_0), .Z(U6_Z_0) );
  IV U194 ( .A(n30), .Z(n426) );
  IV U195 ( .A(n33), .Z(n425) );
  IV U196 ( .A(n46), .Z(n424) );
  IV U197 ( .A(n60), .Z(n423) );
  IV U198 ( .A(n65), .Z(n422) );
  IV U199 ( .A(n69), .Z(n421) );
  IV U200 ( .A(n49), .Z(n419) );
  IV U201 ( .A(n74), .Z(n418) );
  IV U202 ( .A(n76), .Z(n417) );
  IV U203 ( .A(n78), .Z(n416) );
  IV U204 ( .A(n80), .Z(n415) );
  IV U205 ( .A(n82), .Z(n414) );
  IV U206 ( .A(n84), .Z(n413) );
  IV U207 ( .A(n87), .Z(n412) );
  IV U208 ( .A(n52), .Z(n410) );
  IV U209 ( .A(n89), .Z(n409) );
  IV U210 ( .A(n91), .Z(n408) );
  IV U211 ( .A(n94), .Z(n407) );
  IV U212 ( .A(n98), .Z(n406) );
  IV U213 ( .A(n102), .Z(n405) );
  IV U214 ( .A(n106), .Z(n404) );
  IV U215 ( .A(n108), .Z(n403) );
  IV U216 ( .A(n19), .Z(n402) );
  IV U217 ( .A(n26), .Z(n399) );
  IV U218 ( .A(n41), .Z(n398) );
  IV U219 ( .A(n44), .Z(n396) );
  IV U220 ( .A(n195), .Z(n395) );
  IV U221 ( .A(n37), .Z(n392) );
  IV U222 ( .A(n13), .Z(n391) );
  OR2 U223 ( .A(n435), .B(n344), .Z(n390) );
  AN2 U224 ( .A(n327), .B(n196), .Z(n435) );
  OR2 U225 ( .A(n436), .B(n342), .Z(n389) );
  AN2 U226 ( .A(n327), .B(n195), .Z(n436) );
  OR2 U227 ( .A(n437), .B(n340), .Z(n388) );
  AN2 U228 ( .A(n327), .B(n204), .Z(n437) );
  OR2 U229 ( .A(n438), .B(n338), .Z(n387) );
  AN2 U230 ( .A(n327), .B(n203), .Z(n438) );
  OR2 U231 ( .A(n439), .B(n336), .Z(n386) );
  AN2 U232 ( .A(n327), .B(n202), .Z(n439) );
  OR2 U233 ( .A(n440), .B(n334), .Z(n385) );
  AN2 U234 ( .A(n327), .B(n201), .Z(n440) );
  OR2 U235 ( .A(n441), .B(n332), .Z(n384) );
  AN2 U236 ( .A(n327), .B(n200), .Z(n441) );
  OR2 U237 ( .A(n442), .B(n330), .Z(n383) );
  AN2 U238 ( .A(n327), .B(n199), .Z(n442) );
  OR2 U239 ( .A(n443), .B(n328), .Z(n382) );
  AN2 U240 ( .A(n327), .B(n198), .Z(n443) );
  OR2 U241 ( .A(n444), .B(n325), .Z(n381) );
  AN2 U242 ( .A(n327), .B(n197), .Z(n444) );
  OR2 U243 ( .A(n445), .B(n446), .Z(n380) );
  OR2 U244 ( .A(n447), .B(n448), .Z(n446) );
  AN2 U245 ( .A(HSS_TXD[7]), .B(n449), .Z(n448) );
  AN2 U246 ( .A(RX_LoopbackData_P2[7]), .B(n450), .Z(n447) );
  OR2 U247 ( .A(n451), .B(n452), .Z(n445) );
  AN2 U248 ( .A(n453), .B(n15), .Z(n452) );
  AN2 U249 ( .A(n454), .B(n455), .Z(n451) );
  IV U250 ( .A(n15), .Z(n455) );
  OR2 U251 ( .A(n456), .B(n457), .Z(n379) );
  OR2 U252 ( .A(n458), .B(n459), .Z(n457) );
  AN2 U253 ( .A(HSS_TXD[8]), .B(n449), .Z(n459) );
  AN2 U254 ( .A(RX_LoopbackData_P2[8]), .B(n450), .Z(n458) );
  OR2 U255 ( .A(n460), .B(n461), .Z(n456) );
  AN2 U256 ( .A(n453), .B(n204), .Z(n461) );
  AN2 U257 ( .A(n454), .B(n397), .Z(n460) );
  IV U258 ( .A(n204), .Z(n397) );
  OR2 U259 ( .A(n462), .B(n463), .Z(n378) );
  OR2 U260 ( .A(n464), .B(n465), .Z(n463) );
  AN2 U261 ( .A(RX_LoopbackData_P2[4]), .B(n450), .Z(n465) );
  AN2 U262 ( .A(n466), .B(U5_DATA2_4), .Z(n464) );
  AN2 U263 ( .A(HSS_TXD[4]), .B(n449), .Z(n462) );
  OR2 U264 ( .A(n467), .B(n468), .Z(n377) );
  OR2 U265 ( .A(n469), .B(n470), .Z(n468) );
  AN2 U266 ( .A(HSS_TXD[9]), .B(n449), .Z(n470) );
  AN2 U267 ( .A(RX_LoopbackData_P2[9]), .B(n450), .Z(n469) );
  OR2 U268 ( .A(n471), .B(n472), .Z(n467) );
  AN2 U269 ( .A(n16), .B(n453), .Z(n472) );
  AN2 U270 ( .A(n454), .B(n473), .Z(n471) );
  IV U271 ( .A(n16), .Z(n473) );
  OR2 U272 ( .A(n474), .B(n475), .Z(n376) );
  OR2 U273 ( .A(n476), .B(n477), .Z(n475) );
  AN2 U274 ( .A(HSS_TXD[6]), .B(n449), .Z(n477) );
  AN2 U275 ( .A(RX_LoopbackData_P2[6]), .B(n450), .Z(n476) );
  OR2 U276 ( .A(n478), .B(n479), .Z(n474) );
  AN2 U277 ( .A(n14), .B(n453), .Z(n479) );
  AN2 U278 ( .A(n480), .B(n466), .Z(n453) );
  IV U279 ( .A(n22), .Z(n480) );
  AN2 U280 ( .A(n454), .B(n481), .Z(n478) );
  IV U281 ( .A(n14), .Z(n481) );
  AN2 U282 ( .A(n466), .B(n22), .Z(n454) );
  OR2 U283 ( .A(n482), .B(n483), .Z(n375) );
  OR2 U284 ( .A(n484), .B(n485), .Z(n483) );
  AN2 U285 ( .A(RX_LoopbackData_P2[5]), .B(n450), .Z(n485) );
  AN2 U286 ( .A(n466), .B(U5_DATA2_5), .Z(n484) );
  AN2 U287 ( .A(HSS_TXD[5]), .B(n449), .Z(n482) );
  OR2 U288 ( .A(n486), .B(n487), .Z(n374) );
  OR2 U289 ( .A(n488), .B(n489), .Z(n487) );
  AN2 U290 ( .A(HSS_TXD[0]), .B(n449), .Z(n489) );
  AN2 U291 ( .A(RX_LoopbackData_P2[0]), .B(n450), .Z(n488) );
  OR2 U292 ( .A(n490), .B(n491), .Z(n486) );
  AN2 U293 ( .A(n492), .B(n197), .Z(n491) );
  AN2 U294 ( .A(n493), .B(n429), .Z(n490) );
  OR2 U295 ( .A(n494), .B(n495), .Z(n373) );
  OR2 U296 ( .A(n496), .B(n497), .Z(n495) );
  AN2 U297 ( .A(HSS_TXD[1]), .B(n449), .Z(n497) );
  AN2 U298 ( .A(RX_LoopbackData_P2[1]), .B(n450), .Z(n496) );
  OR2 U299 ( .A(n498), .B(n499), .Z(n494) );
  AN2 U300 ( .A(n[5]), .B(n492), .Z(n499) );
  AN2 U301 ( .A(n493), .B(n500), .Z(n498) );
  IV U302 ( .A(n[5]), .Z(n500) );
  OR2 U303 ( .A(n501), .B(n502), .Z(n372) );
  OR2 U304 ( .A(n503), .B(n504), .Z(n502) );
  AN2 U305 ( .A(HSS_TXD[2]), .B(n449), .Z(n504) );
  AN2 U306 ( .A(RX_LoopbackData_P2[2]), .B(n450), .Z(n503) );
  OR2 U307 ( .A(n505), .B(n506), .Z(n501) );
  AN2 U308 ( .A(n[6]), .B(n492), .Z(n506) );
  AN2 U309 ( .A(n493), .B(n507), .Z(n505) );
  IV U310 ( .A(n[6]), .Z(n507) );
  OR2 U311 ( .A(n508), .B(n509), .Z(n371) );
  OR2 U312 ( .A(n510), .B(n511), .Z(n509) );
  AN2 U313 ( .A(HSS_TXD[3]), .B(n449), .Z(n511) );
  AN2 U314 ( .A(RX_LoopbackData_P2[3]), .B(n450), .Z(n510) );
  AN2 U315 ( .A(n194), .B(CNTL_Loopback_P0), .Z(n450) );
  OR2 U316 ( .A(n512), .B(n513), .Z(n508) );
  AN2 U317 ( .A(n[7]), .B(n492), .Z(n513) );
  AN2 U318 ( .A(n514), .B(n466), .Z(n492) );
  AN2 U319 ( .A(n493), .B(n515), .Z(n512) );
  IV U320 ( .A(n[7]), .Z(n515) );
  AN2 U321 ( .A(n466), .B(n21), .Z(n493) );
  AN2 U322 ( .A(n181), .B(n194), .Z(n466) );
  OR2 U323 ( .A(n516), .B(n517), .Z(n154) );
  IV U324 ( .A(n518), .Z(n517) );
  OR2 U325 ( .A(n434), .B(n153), .Z(n518) );
  AN2 U326 ( .A(n153), .B(n434), .Z(n516) );
  IV U327 ( .A(n393), .Z(n434) );
  OR2 U328 ( .A(n519), .B(n520), .Z(n393) );
  AN2 U329 ( .A(n151), .B(n394), .Z(n520) );
  IV U330 ( .A(n521), .Z(n519) );
  OR2 U331 ( .A(n394), .B(n151), .Z(n521) );
  IV U332 ( .A(n20), .Z(n394) );
  OR2 U333 ( .A(n522), .B(n523), .Z(n147) );
  AN2 U334 ( .A(n202), .B(n400), .Z(n523) );
  IV U335 ( .A(n203), .Z(n400) );
  AN2 U336 ( .A(n203), .B(n401), .Z(n522) );
  IV U337 ( .A(n202), .Z(n401) );
  OR2 U338 ( .A(n524), .B(n525), .Z(n119) );
  AN2 U339 ( .A(n199), .B(n420), .Z(n525) );
  IV U340 ( .A(n200), .Z(n420) );
  AN2 U341 ( .A(n200), .B(n427), .Z(n524) );
  IV U342 ( .A(n199), .Z(n427) );
  OR2 U343 ( .A(n526), .B(n527), .Z(n118) );
  AN2 U344 ( .A(n197), .B(n428), .Z(n527) );
  IV U345 ( .A(n198), .Z(n428) );
  AN2 U346 ( .A(n198), .B(n429), .Z(n526) );
  IV U347 ( .A(n197), .Z(n429) );
  OR2 U348 ( .A(n528), .B(n529), .Z(n116) );
  IV U349 ( .A(n530), .Z(n529) );
  OR2 U350 ( .A(n411), .B(n28), .Z(n530) );
  AN2 U351 ( .A(n28), .B(n411), .Z(n528) );
  AN2 U352 ( .A(n531), .B(n532), .Z(n113) );
  IV U353 ( .A(n533), .Z(n532) );
  AN2 U354 ( .A(n411), .B(n55), .Z(n533) );
  OR2 U355 ( .A(n55), .B(n411), .Z(n531) );
  IV U356 ( .A(n201), .Z(n411) );
  OR2 U357 ( .A(n534), .B(n535), .Z(U5_DATA2_5) );
  IV U358 ( .A(n536), .Z(n535) );
  OR2 U359 ( .A(n514), .B(n[9]), .Z(n536) );
  AN2 U360 ( .A(n[9]), .B(n514), .Z(n534) );
  OR2 U361 ( .A(n537), .B(n538), .Z(U5_DATA2_4) );
  IV U362 ( .A(n539), .Z(n538) );
  OR2 U363 ( .A(n514), .B(n[8]), .Z(n539) );
  AN2 U364 ( .A(n[8]), .B(n514), .Z(n537) );
  IV U365 ( .A(n21), .Z(n514) );
  OR2 U366 ( .A(n540), .B(n168), .Z(U4_Z_0) );
  AN2 U367 ( .A(CNTL_RESETN_P0), .B(n449), .Z(n540) );
  IV U368 ( .A(n194), .Z(n449) );
endmodule

