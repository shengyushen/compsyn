
module PCIEXP_TX ( PCLK250, RST_BeaconEnable_R0, CNTL_RESETN_P0, 
        CNTL_Loopback_P0, CNTL_TXEnable_P0, RX_LoopbackData_P2, TXCOMPLIANCE, 
        TXDATA, TXDATAK, TXELECIDLE, HSS_TXBEACONCMD, HSS_TXD, HSS_TXELECIDLE, 
        assertion_shengyushen );
  input [9:0] RX_LoopbackData_P2;
  input [7:0] TXDATA;
  output [9:0] HSS_TXD;
  input PCLK250, RST_BeaconEnable_R0, CNTL_RESETN_P0, CNTL_Loopback_P0,
         CNTL_TXEnable_P0, TXCOMPLIANCE, TXDATAK, TXELECIDLE;
  output HSS_TXBEACONCMD, HSS_TXELECIDLE, assertion_shengyushen;
  wire   n3, n4, n10, n11, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n25, n26, n28, n29, n30, n31, n32, n33, n35, n36, n37, n39, n40, n41,
         n44, n46, n48, n49, n52, n55, n58, n59, n60, n63, n64, n65, n68, n69,
         n71, n72, n73, n74, n76, n78, n80, n82, n84, n86, n87, n89, n91, n93,
         n94, n96, n97, n98, n100, n101, n102, n104, n105, n106, n108, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n140, n141, n142, n145, n146, n147,
         n148, n149, n150, n151, n153, n154, n157, n158, n159, n160, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n280, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, U6_Z_0, U6_DATA2_0,
         U5_DATA2_4, U5_DATA2_5, U4_Z_0, n425, n427, n428, n430, n432, n434,
         n436, n438, n440, n442, n444, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640;
  wire   [5:9] n;

  OR2 C36 ( .A(n500), .B(n501), .Z(n25) );
  OR2 C37 ( .A(n303), .B(n25), .Z(n26) );
  AN2 C39 ( .A(n297), .B(n296), .Z(n28) );
  AN2 C40 ( .A(n298), .B(n28), .Z(n29) );
  AN2 C41 ( .A(n299), .B(n29), .Z(n30) );
  OR2 C42 ( .A(n297), .B(n296), .Z(n31) );
  OR2 C43 ( .A(n298), .B(n31), .Z(n32) );
  OR2 C44 ( .A(n299), .B(n32), .Z(n33) );
  AN2 C46 ( .A(n302), .B(n301), .Z(n35) );
  AN2 C47 ( .A(n303), .B(n35), .Z(n36) );
  OR2 C48 ( .A(U5_DATA2_5), .B(U5_DATA2_4), .Z(n37) );
  AN2 C50 ( .A(U5_DATA2_5), .B(U5_DATA2_4), .Z(n39) );
  OR2 C53 ( .A(n302), .B(n301), .Z(n40) );
  OR2 C54 ( .A(n303), .B(n40), .Z(n41) );
  OR2 C58 ( .A(n497), .B(n40), .Z(n44) );
  OR2 C60 ( .A(n299), .B(n298), .Z(n46) );
  OR2 C67 ( .A(n520), .B(n68), .Z(n48) );
  OR2 C68 ( .A(n300), .B(n48), .Z(n49) );
  OR2 C75 ( .A(n511), .B(n69), .Z(n52) );
  OR2 C80 ( .A(n520), .B(n32), .Z(n55) );
  OR2 C83 ( .A(n297), .B(n529), .Z(n58) );
  OR2 C84 ( .A(n298), .B(n58), .Z(n59) );
  OR2 C85 ( .A(n299), .B(n59), .Z(n60) );
  OR2 C88 ( .A(n528), .B(n296), .Z(n63) );
  OR2 C89 ( .A(n298), .B(n63), .Z(n64) );
  OR2 C90 ( .A(n299), .B(n64), .Z(n65) );
  OR2 C941 ( .A(n527), .B(n31), .Z(n68) );
  OR2 C951 ( .A(n299), .B(n68), .Z(n69) );
  OR2 C100 ( .A(n528), .B(n529), .Z(n71) );
  OR2 C101 ( .A(n527), .B(n71), .Z(n72) );
  OR2 C102 ( .A(n299), .B(n72), .Z(n73) );
  OR2 C103 ( .A(n300), .B(n73), .Z(n74) );
  OR2 C1081 ( .A(n300), .B(n33), .Z(n76) );
  OR2 C114 ( .A(n300), .B(n60), .Z(n78) );
  OR2 C1201 ( .A(n300), .B(n65), .Z(n80) );
  OR2 C126 ( .A(n300), .B(n69), .Z(n82) );
  OR2 C1321 ( .A(n300), .B(n55), .Z(n84) );
  OR2 C140 ( .A(n520), .B(n72), .Z(n86) );
  OR2 C141 ( .A(n300), .B(n86), .Z(n87) );
  OR2 C1481 ( .A(n511), .B(n55), .Z(n89) );
  OR2 C154 ( .A(n511), .B(n33), .Z(n91) );
  AN2 C1591 ( .A(n300), .B(n30), .Z(n93) );
  OR2 C167 ( .A(n511), .B(n73), .Z(n94) );
  OR2 C1741 ( .A(n298), .B(n71), .Z(n96) );
  OR2 C175 ( .A(n520), .B(n96), .Z(n97) );
  OR2 C176 ( .A(n511), .B(n97), .Z(n98) );
  OR2 C1831 ( .A(n527), .B(n58), .Z(n100) );
  OR2 C1841 ( .A(n520), .B(n100), .Z(n101) );
  OR2 C1851 ( .A(n511), .B(n101), .Z(n102) );
  OR2 C192 ( .A(n527), .B(n63), .Z(n104) );
  OR2 C193 ( .A(n520), .B(n104), .Z(n105) );
  OR2 C194 ( .A(n511), .B(n105), .Z(n106) );
  OR2 C2021 ( .A(n511), .B(n48), .Z(n108) );
  OR2 C206 ( .A(n111), .B(n525), .Z(n[5]) );
  AN2 C207 ( .A(n297), .B(n526), .Z(n111) );
  OR2 C209 ( .A(n112), .B(n509), .Z(n[6]) );
  OR2 C210 ( .A(n298), .B(n525), .Z(n112) );
  AN2 C211 ( .A(n299), .B(n526), .Z(n[7]) );
  OR2 C213 ( .A(n113), .B(n115), .Z(n[8]) );
  OR2 C215 ( .A(n114), .B(n521), .Z(n115) );
  OR2 C2161 ( .A(n523), .B(n522), .Z(n114) );
  OR2 C2171 ( .A(n125), .B(n126), .Z(n[9]) );
  OR2 C2181 ( .A(n124), .B(n93), .Z(n125) );
  OR2 C219 ( .A(n123), .B(n510), .Z(n124) );
  OR2 C220 ( .A(n122), .B(n519), .Z(n123) );
  OR2 C221 ( .A(n117), .B(n121), .Z(n122) );
  AN2 C222 ( .A(n524), .B(n116), .Z(n117) );
  AN2 C224 ( .A(n120), .B(n511), .Z(n121) );
  AN2 C225 ( .A(n118), .B(n119), .Z(n120) );
  AN2 C229 ( .A(n503), .B(n295), .Z(n126) );
  OR2 C230 ( .A(n131), .B(n509), .Z(n10) );
  OR2 C231 ( .A(n130), .B(n512), .Z(n131) );
  OR2 C232 ( .A(n129), .B(n513), .Z(n130) );
  OR2 C2331 ( .A(n128), .B(n514), .Z(n129) );
  OR2 C234 ( .A(n127), .B(n515), .Z(n128) );
  OR2 C235 ( .A(n517), .B(n516), .Z(n127) );
  OR2 C236 ( .A(n136), .B(n137), .Z(n11) );
  OR2 C237 ( .A(n135), .B(n93), .Z(n136) );
  OR2 C238 ( .A(n134), .B(n504), .Z(n135) );
  OR2 C239 ( .A(n133), .B(n505), .Z(n134) );
  OR2 C240 ( .A(n132), .B(n506), .Z(n133) );
  OR2 C241 ( .A(n508), .B(n507), .Z(n132) );
  AN2 C242 ( .A(n503), .B(n295), .Z(n137) );
  AN2 C243 ( .A(n142), .B(n36), .Z(n13) );
  OR2 C244 ( .A(n141), .B(n295), .Z(n142) );
  OR2 C245 ( .A(n138), .B(n140), .Z(n141) );
  AN2 C246 ( .A(n493), .B(n492), .Z(n138) );
  AN2 C2471 ( .A(n534), .B(n39), .Z(n140) );
  AN2 C249 ( .A(n301), .B(n491), .Z(n14) );
  OR2 C251 ( .A(n302), .B(n498), .Z(n15) );
  OR2 C2521 ( .A(n145), .B(n13), .Z(n16) );
  AN2 C2531 ( .A(n147), .B(n497), .Z(n145) );
  OR2 C256 ( .A(n498), .B(n496), .Z(n17) );
  AN2 C2571 ( .A(n146), .B(n147), .Z(n18) );
  AN2 C258 ( .A(n503), .B(n295), .Z(n146) );
  OR2 C260 ( .A(n150), .B(n503), .Z(n19) );
  OR2 C261 ( .A(n149), .B(n504), .Z(n150) );
  OR2 C262 ( .A(n148), .B(n505), .Z(n149) );
  OR2 C263 ( .A(n507), .B(n506), .Z(n148) );
  OR2 C265 ( .A(n10), .B(n11), .Z(n151) );
  AN2 C266 ( .A(n293), .B(n154), .Z(n4) );
  OR2 C269 ( .A(n17), .B(n36), .Z(n153) );
  AN2 C2701 ( .A(n495), .B(n3), .Z(n20) );
  OR2 C2721 ( .A(n160), .B(n162), .Z(n21) );
  OR2 C2731 ( .A(n157), .B(n159), .Z(n160) );
  AN2 C2741 ( .A(n494), .B(n10), .Z(n157) );
  AN2 C2761 ( .A(n20), .B(n158), .Z(n159) );
  OR2 C2771 ( .A(n518), .B(n11), .Z(n158) );
  AN2 C2781 ( .A(n502), .B(n295), .Z(n162) );
  OR2 C2801 ( .A(n164), .B(n166), .Z(n22) );
  AN2 C2811 ( .A(n534), .B(n163), .Z(n164) );
  OR2 C2831 ( .A(n17), .B(n18), .Z(n163) );
  AN2 C2841 ( .A(n493), .B(n165), .Z(n166) );
  OR2 C2851 ( .A(n499), .B(n36), .Z(n165) );
  OR2 C286 ( .A(n256), .B(n248), .Z(n182) );
  OR2 C285 ( .A(n182), .B(n239), .Z(n181) );
  OR2 C284 ( .A(n181), .B(n232), .Z(n180) );
  OR2 C283 ( .A(n180), .B(n223), .Z(n179) );
  OR2 C282 ( .A(n179), .B(n216), .Z(n178) );
  OR2 C281 ( .A(n178), .B(n208), .Z(n177) );
  OR2 C280 ( .A(n177), .B(n201), .Z(n176) );
  OR2 C279 ( .A(n176), .B(n194), .Z(n175) );
  OR2 C278 ( .A(n175), .B(n190), .Z(n174) );
  OR2 C277 ( .A(n174), .B(n188), .Z(n173) );
  OR2 C276 ( .A(n173), .B(n185), .Z(n172) );
  AN2 C275 ( .A(TXDATAK), .B(n172), .Z(n171) );
  OR2 C274 ( .A(n267), .B(n171), .Z(n170) );
  AN2 C273 ( .A(n170), .B(CNTL_RESETN_P0), .Z(n169) );
  AN2 C272 ( .A(n169), .B(n280), .Z(n168) );
  AN2 C271 ( .A(n168), .B(n183), .Z(n167) );
  AN2 C270 ( .A(n167), .B(CNTL_TXEnable_P0), .Z(assertion_shengyushen) );
  IV I_24 ( .A(CNTL_Loopback_P0), .Z(n280) );
  AN2 C259 ( .A(CNTL_TXEnable_P0), .B(n183), .Z(U6_DATA2_0) );
  IV I_22 ( .A(TXELECIDLE), .Z(n183) );
  AN2 C257 ( .A(RST_BeaconEnable_R0), .B(n183), .Z(HSS_TXBEACONCMD) );
  IV I_21 ( .A(CNTL_RESETN_P0), .Z(n184) );
  IV I_20 ( .A(n186), .Z(n185) );
  OR2 C248 ( .A(TXDATA[0]), .B(n187), .Z(n186) );
  OR2 C247 ( .A(n200), .B(n204), .Z(n187) );
  IV I_19 ( .A(n189), .Z(n188) );
  OR2 C233 ( .A(n199), .B(n203), .Z(n189) );
  IV I_18 ( .A(n191), .Z(n190) );
  OR2 C218 ( .A(n199), .B(n192), .Z(n191) );
  OR2 C217 ( .A(n200), .B(n193), .Z(n192) );
  OR2 C216 ( .A(TXDATA[2]), .B(n205), .Z(n193) );
  IV I_17 ( .A(n195), .Z(n194) );
  OR2 C203 ( .A(n199), .B(n196), .Z(n195) );
  OR2 C202 ( .A(n200), .B(n197), .Z(n196) );
  OR2 C201 ( .A(n264), .B(n198), .Z(n197) );
  OR2 C200 ( .A(TXDATA[3]), .B(n206), .Z(n198) );
  IV I_16 ( .A(TXDATA[0]), .Z(n199) );
  IV I_15 ( .A(TXDATA[1]), .Z(n200) );
  IV I_14 ( .A(n202), .Z(n201) );
  OR2 C188 ( .A(TXDATA[0]), .B(n203), .Z(n202) );
  OR2 C187 ( .A(TXDATA[1]), .B(n204), .Z(n203) );
  OR2 C186 ( .A(n264), .B(n205), .Z(n204) );
  OR2 C185 ( .A(n265), .B(n206), .Z(n205) );
  OR2 C184 ( .A(n266), .B(n207), .Z(n206) );
  OR2 C183 ( .A(n255), .B(n215), .Z(n207) );
  IV I_13 ( .A(n209), .Z(n208) );
  OR2 C174 ( .A(TXDATA[0]), .B(n210), .Z(n209) );
  OR2 C173 ( .A(TXDATA[1]), .B(n211), .Z(n210) );
  OR2 C172 ( .A(n264), .B(n212), .Z(n211) );
  OR2 C171 ( .A(n265), .B(n213), .Z(n212) );
  OR2 C170 ( .A(n266), .B(n214), .Z(n213) );
  OR2 C169 ( .A(TXDATA[5]), .B(n215), .Z(n214) );
  OR2 C168 ( .A(n247), .B(n231), .Z(n215) );
  IV I_12 ( .A(n217), .Z(n216) );
  OR2 C161 ( .A(TXDATA[0]), .B(n218), .Z(n217) );
  OR2 C160 ( .A(TXDATA[1]), .B(n219), .Z(n218) );
  OR2 C159 ( .A(n264), .B(n220), .Z(n219) );
  OR2 C158 ( .A(n265), .B(n221), .Z(n220) );
  OR2 C157 ( .A(n266), .B(n222), .Z(n221) );
  OR2 C156 ( .A(n255), .B(n230), .Z(n222) );
  IV I_11 ( .A(n224), .Z(n223) );
  OR2 C148 ( .A(TXDATA[0]), .B(n225), .Z(n224) );
  OR2 C147 ( .A(TXDATA[1]), .B(n226), .Z(n225) );
  OR2 C146 ( .A(n264), .B(n227), .Z(n226) );
  OR2 C145 ( .A(n265), .B(n228), .Z(n227) );
  OR2 C144 ( .A(n266), .B(n229), .Z(n228) );
  OR2 C143 ( .A(TXDATA[5]), .B(n230), .Z(n229) );
  OR2 C142 ( .A(TXDATA[6]), .B(n231), .Z(n230) );
  IV I_10 ( .A(TXDATA[7]), .Z(n231) );
  IV I_9 ( .A(n233), .Z(n232) );
  OR2 C136 ( .A(TXDATA[0]), .B(n234), .Z(n233) );
  OR2 C135 ( .A(TXDATA[1]), .B(n235), .Z(n234) );
  OR2 C134 ( .A(n264), .B(n236), .Z(n235) );
  OR2 C133 ( .A(n265), .B(n237), .Z(n236) );
  OR2 C132 ( .A(n266), .B(n238), .Z(n237) );
  OR2 C131 ( .A(n255), .B(n246), .Z(n238) );
  IV I_8 ( .A(n240), .Z(n239) );
  OR2 C123 ( .A(TXDATA[0]), .B(n241), .Z(n240) );
  OR2 C122 ( .A(TXDATA[1]), .B(n242), .Z(n241) );
  OR2 C121 ( .A(n264), .B(n243), .Z(n242) );
  OR2 C120 ( .A(n265), .B(n244), .Z(n243) );
  OR2 C119 ( .A(n266), .B(n245), .Z(n244) );
  OR2 C118 ( .A(TXDATA[5]), .B(n246), .Z(n245) );
  OR2 C117 ( .A(n247), .B(TXDATA[7]), .Z(n246) );
  IV I_7 ( .A(TXDATA[6]), .Z(n247) );
  IV I_6 ( .A(n249), .Z(n248) );
  OR2 C111 ( .A(TXDATA[0]), .B(n250), .Z(n249) );
  OR2 C110 ( .A(TXDATA[1]), .B(n251), .Z(n250) );
  OR2 C109 ( .A(n264), .B(n252), .Z(n251) );
  OR2 C108 ( .A(n265), .B(n253), .Z(n252) );
  OR2 C107 ( .A(n266), .B(n254), .Z(n253) );
  OR2 C106 ( .A(n255), .B(n263), .Z(n254) );
  IV I_5 ( .A(TXDATA[5]), .Z(n255) );
  IV I_4 ( .A(n257), .Z(n256) );
  OR2 C99 ( .A(TXDATA[0]), .B(n258), .Z(n257) );
  OR2 C98 ( .A(TXDATA[1]), .B(n259), .Z(n258) );
  OR2 C97 ( .A(n264), .B(n260), .Z(n259) );
  OR2 C96 ( .A(n265), .B(n261), .Z(n260) );
  OR2 C95 ( .A(n266), .B(n262), .Z(n261) );
  OR2 C94 ( .A(TXDATA[5]), .B(n263), .Z(n262) );
  OR2 C93 ( .A(TXDATA[6]), .B(TXDATA[7]), .Z(n263) );
  IV I_3 ( .A(TXDATA[2]), .Z(n264) );
  IV I_2 ( .A(TXDATA[3]), .Z(n265) );
  IV I_1 ( .A(TXDATA[4]), .Z(n266) );
  IV I_0 ( .A(TXDATAK), .Z(n267) );
  FD1 InputDataK_P0_reg ( .D(n490), .CP(PCLK250), .Q(n295) );
  FD1 InputCompliance_P0_reg ( .D(n489), .CP(PCLK250), .Q(n294) );
  FD1 InputData_P0_reg_7_ ( .D(n488), .CP(PCLK250), .Q(n303) );
  FD1 InputData_P0_reg_6_ ( .D(n487), .CP(PCLK250), .Q(n302) );
  FD1 InputData_P0_reg_5_ ( .D(n486), .CP(PCLK250), .Q(n301) );
  FD1 InputData_P0_reg_4_ ( .D(n485), .CP(PCLK250), .Q(n300) );
  FD1 InputData_P0_reg_3_ ( .D(n484), .CP(PCLK250), .Q(n299) );
  FD1 InputData_P0_reg_2_ ( .D(n483), .CP(PCLK250), .Q(n298) );
  FD1 InputData_P0_reg_1_ ( .D(n482), .CP(PCLK250), .Q(n297) );
  FD1 InputData_P0_reg_0_ ( .D(n481), .CP(PCLK250), .Q(n296) );
  FD1 InputDataEnable_P0_reg ( .D(U6_Z_0), .CP(PCLK250), .Q(n293) );
  FD1 OutputElecIdle_P0_reg ( .D(U4_Z_0), .CP(PCLK250), .Q(HSS_TXELECIDLE) );
  FD1 DISPARITY_P0_reg ( .D(n4), .CP(PCLK250), .Q(n3) );
  FD1 OutputData_P0_reg_7_ ( .D(n480), .CP(PCLK250), .Q(HSS_TXD[7]) );
  FD1 OutputData_P0_reg_8_ ( .D(n479), .CP(PCLK250), .Q(HSS_TXD[8]) );
  FD1 OutputData_P0_reg_4_ ( .D(n478), .CP(PCLK250), .Q(HSS_TXD[4]) );
  FD1 OutputData_P0_reg_9_ ( .D(n477), .CP(PCLK250), .Q(HSS_TXD[9]) );
  FD1 OutputData_P0_reg_6_ ( .D(n476), .CP(PCLK250), .Q(HSS_TXD[6]) );
  FD1 OutputData_P0_reg_5_ ( .D(n475), .CP(PCLK250), .Q(HSS_TXD[5]) );
  FD1 OutputData_P0_reg_0_ ( .D(n474), .CP(PCLK250), .Q(HSS_TXD[0]) );
  FD1 OutputData_P0_reg_1_ ( .D(n473), .CP(PCLK250), .Q(HSS_TXD[1]) );
  FD1 OutputData_P0_reg_2_ ( .D(n472), .CP(PCLK250), .Q(HSS_TXD[2]) );
  FD1 OutputData_P0_reg_3_ ( .D(n471), .CP(PCLK250), .Q(HSS_TXD[3]) );
  AN2 U88 ( .A(U6_DATA2_0), .B(TXDATA[0]), .Z(n425) );
  AN2 U91 ( .A(TXDATA[1]), .B(U6_DATA2_0), .Z(n428) );
  AN2 U94 ( .A(TXDATA[2]), .B(U6_DATA2_0), .Z(n430) );
  AN2 U97 ( .A(TXDATA[3]), .B(U6_DATA2_0), .Z(n432) );
  AN2 U100 ( .A(TXDATA[4]), .B(U6_DATA2_0), .Z(n434) );
  AN2 U103 ( .A(TXDATA[5]), .B(U6_DATA2_0), .Z(n436) );
  AN2 U106 ( .A(TXDATA[6]), .B(U6_DATA2_0), .Z(n438) );
  AN2 U109 ( .A(TXDATA[7]), .B(U6_DATA2_0), .Z(n440) );
  AN2 U112 ( .A(TXCOMPLIANCE), .B(U6_DATA2_0), .Z(n442) );
  IV U115 ( .A(U6_DATA2_0), .Z(n427) );
  AN2 U116 ( .A(TXDATAK), .B(U6_DATA2_0), .Z(n444) );
  AN2 U181 ( .A(CNTL_RESETN_P0), .B(U6_DATA2_0), .Z(U6_Z_0) );
  IV U194 ( .A(n30), .Z(n526) );
  IV U195 ( .A(n33), .Z(n525) );
  IV U196 ( .A(n46), .Z(n524) );
  IV U197 ( .A(n60), .Z(n523) );
  IV U198 ( .A(n65), .Z(n522) );
  IV U199 ( .A(n69), .Z(n521) );
  IV U200 ( .A(n49), .Z(n519) );
  IV U201 ( .A(n74), .Z(n518) );
  IV U202 ( .A(n76), .Z(n517) );
  IV U203 ( .A(n78), .Z(n516) );
  IV U204 ( .A(n80), .Z(n515) );
  IV U205 ( .A(n82), .Z(n514) );
  IV U206 ( .A(n84), .Z(n513) );
  IV U207 ( .A(n87), .Z(n512) );
  IV U208 ( .A(n52), .Z(n510) );
  IV U209 ( .A(n89), .Z(n509) );
  IV U210 ( .A(n91), .Z(n508) );
  IV U211 ( .A(n94), .Z(n507) );
  IV U212 ( .A(n98), .Z(n506) );
  IV U213 ( .A(n102), .Z(n505) );
  IV U214 ( .A(n106), .Z(n504) );
  IV U215 ( .A(n108), .Z(n503) );
  IV U216 ( .A(n19), .Z(n502) );
  IV U217 ( .A(n26), .Z(n499) );
  IV U218 ( .A(n41), .Z(n498) );
  IV U219 ( .A(n44), .Z(n496) );
  IV U220 ( .A(n294), .Z(n495) );
  IV U221 ( .A(n37), .Z(n492) );
  IV U222 ( .A(n13), .Z(n491) );
  OR2 U223 ( .A(n535), .B(n444), .Z(n490) );
  AN2 U224 ( .A(n427), .B(n295), .Z(n535) );
  OR2 U225 ( .A(n536), .B(n442), .Z(n489) );
  AN2 U226 ( .A(n427), .B(n294), .Z(n536) );
  OR2 U227 ( .A(n537), .B(n440), .Z(n488) );
  AN2 U228 ( .A(n427), .B(n303), .Z(n537) );
  OR2 U229 ( .A(n538), .B(n438), .Z(n487) );
  AN2 U230 ( .A(n427), .B(n302), .Z(n538) );
  OR2 U231 ( .A(n539), .B(n436), .Z(n486) );
  AN2 U232 ( .A(n427), .B(n301), .Z(n539) );
  OR2 U233 ( .A(n540), .B(n434), .Z(n485) );
  AN2 U234 ( .A(n427), .B(n300), .Z(n540) );
  OR2 U235 ( .A(n541), .B(n432), .Z(n484) );
  AN2 U236 ( .A(n427), .B(n299), .Z(n541) );
  OR2 U237 ( .A(n542), .B(n430), .Z(n483) );
  AN2 U238 ( .A(n427), .B(n298), .Z(n542) );
  OR2 U239 ( .A(n543), .B(n428), .Z(n482) );
  AN2 U240 ( .A(n427), .B(n297), .Z(n543) );
  OR2 U241 ( .A(n544), .B(n425), .Z(n481) );
  AN2 U242 ( .A(n427), .B(n296), .Z(n544) );
  OR2 U243 ( .A(n545), .B(n546), .Z(n480) );
  OR2 U244 ( .A(n547), .B(n548), .Z(n546) );
  AN2 U245 ( .A(HSS_TXD[7]), .B(n549), .Z(n548) );
  AN2 U246 ( .A(RX_LoopbackData_P2[7]), .B(n550), .Z(n547) );
  OR2 U247 ( .A(n551), .B(n552), .Z(n545) );
  AN2 U248 ( .A(n553), .B(n15), .Z(n552) );
  AN2 U249 ( .A(n554), .B(n555), .Z(n551) );
  IV U250 ( .A(n15), .Z(n555) );
  OR2 U251 ( .A(n556), .B(n557), .Z(n479) );
  OR2 U252 ( .A(n558), .B(n559), .Z(n557) );
  AN2 U253 ( .A(HSS_TXD[8]), .B(n549), .Z(n559) );
  AN2 U254 ( .A(RX_LoopbackData_P2[8]), .B(n550), .Z(n558) );
  OR2 U255 ( .A(n560), .B(n561), .Z(n556) );
  AN2 U256 ( .A(n553), .B(n303), .Z(n561) );
  AN2 U257 ( .A(n554), .B(n497), .Z(n560) );
  IV U258 ( .A(n303), .Z(n497) );
  OR2 U259 ( .A(n562), .B(n563), .Z(n478) );
  OR2 U260 ( .A(n564), .B(n565), .Z(n563) );
  AN2 U261 ( .A(RX_LoopbackData_P2[4]), .B(n550), .Z(n565) );
  AN2 U262 ( .A(n566), .B(U5_DATA2_4), .Z(n564) );
  AN2 U263 ( .A(HSS_TXD[4]), .B(n549), .Z(n562) );
  OR2 U264 ( .A(n567), .B(n568), .Z(n477) );
  OR2 U265 ( .A(n569), .B(n570), .Z(n568) );
  AN2 U266 ( .A(HSS_TXD[9]), .B(n549), .Z(n570) );
  AN2 U267 ( .A(RX_LoopbackData_P2[9]), .B(n550), .Z(n569) );
  OR2 U268 ( .A(n571), .B(n572), .Z(n567) );
  AN2 U269 ( .A(n16), .B(n553), .Z(n572) );
  AN2 U270 ( .A(n554), .B(n573), .Z(n571) );
  IV U271 ( .A(n16), .Z(n573) );
  OR2 U272 ( .A(n574), .B(n575), .Z(n476) );
  OR2 U273 ( .A(n576), .B(n577), .Z(n575) );
  AN2 U274 ( .A(HSS_TXD[6]), .B(n549), .Z(n577) );
  AN2 U275 ( .A(RX_LoopbackData_P2[6]), .B(n550), .Z(n576) );
  OR2 U276 ( .A(n578), .B(n579), .Z(n574) );
  AN2 U277 ( .A(n14), .B(n553), .Z(n579) );
  AN2 U278 ( .A(n580), .B(n566), .Z(n553) );
  IV U279 ( .A(n22), .Z(n580) );
  AN2 U280 ( .A(n554), .B(n581), .Z(n578) );
  IV U281 ( .A(n14), .Z(n581) );
  AN2 U282 ( .A(n566), .B(n22), .Z(n554) );
  OR2 U283 ( .A(n582), .B(n583), .Z(n475) );
  OR2 U284 ( .A(n584), .B(n585), .Z(n583) );
  AN2 U285 ( .A(RX_LoopbackData_P2[5]), .B(n550), .Z(n585) );
  AN2 U286 ( .A(n566), .B(U5_DATA2_5), .Z(n584) );
  AN2 U287 ( .A(HSS_TXD[5]), .B(n549), .Z(n582) );
  OR2 U288 ( .A(n586), .B(n587), .Z(n474) );
  OR2 U289 ( .A(n588), .B(n589), .Z(n587) );
  AN2 U290 ( .A(HSS_TXD[0]), .B(n549), .Z(n589) );
  AN2 U291 ( .A(RX_LoopbackData_P2[0]), .B(n550), .Z(n588) );
  OR2 U292 ( .A(n590), .B(n591), .Z(n586) );
  AN2 U293 ( .A(n592), .B(n296), .Z(n591) );
  AN2 U294 ( .A(n593), .B(n529), .Z(n590) );
  OR2 U295 ( .A(n594), .B(n595), .Z(n473) );
  OR2 U296 ( .A(n596), .B(n597), .Z(n595) );
  AN2 U297 ( .A(HSS_TXD[1]), .B(n549), .Z(n597) );
  AN2 U298 ( .A(RX_LoopbackData_P2[1]), .B(n550), .Z(n596) );
  OR2 U299 ( .A(n598), .B(n599), .Z(n594) );
  AN2 U300 ( .A(n[5]), .B(n592), .Z(n599) );
  AN2 U301 ( .A(n593), .B(n600), .Z(n598) );
  IV U302 ( .A(n[5]), .Z(n600) );
  OR2 U303 ( .A(n601), .B(n602), .Z(n472) );
  OR2 U304 ( .A(n603), .B(n604), .Z(n602) );
  AN2 U305 ( .A(HSS_TXD[2]), .B(n549), .Z(n604) );
  AN2 U306 ( .A(RX_LoopbackData_P2[2]), .B(n550), .Z(n603) );
  OR2 U307 ( .A(n605), .B(n606), .Z(n601) );
  AN2 U308 ( .A(n[6]), .B(n592), .Z(n606) );
  AN2 U309 ( .A(n593), .B(n607), .Z(n605) );
  IV U310 ( .A(n[6]), .Z(n607) );
  OR2 U311 ( .A(n608), .B(n609), .Z(n471) );
  OR2 U312 ( .A(n610), .B(n611), .Z(n609) );
  AN2 U313 ( .A(HSS_TXD[3]), .B(n549), .Z(n611) );
  AN2 U314 ( .A(RX_LoopbackData_P2[3]), .B(n550), .Z(n610) );
  AN2 U315 ( .A(n293), .B(CNTL_Loopback_P0), .Z(n550) );
  OR2 U316 ( .A(n612), .B(n613), .Z(n608) );
  AN2 U317 ( .A(n[7]), .B(n592), .Z(n613) );
  AN2 U318 ( .A(n614), .B(n566), .Z(n592) );
  AN2 U319 ( .A(n593), .B(n615), .Z(n612) );
  IV U320 ( .A(n[7]), .Z(n615) );
  AN2 U321 ( .A(n566), .B(n21), .Z(n593) );
  AN2 U322 ( .A(n280), .B(n293), .Z(n566) );
  OR2 U323 ( .A(n616), .B(n617), .Z(n154) );
  IV U324 ( .A(n618), .Z(n617) );
  OR2 U325 ( .A(n534), .B(n153), .Z(n618) );
  AN2 U326 ( .A(n153), .B(n534), .Z(n616) );
  IV U327 ( .A(n493), .Z(n534) );
  OR2 U328 ( .A(n619), .B(n620), .Z(n493) );
  AN2 U329 ( .A(n151), .B(n494), .Z(n620) );
  IV U330 ( .A(n621), .Z(n619) );
  OR2 U331 ( .A(n494), .B(n151), .Z(n621) );
  IV U332 ( .A(n20), .Z(n494) );
  OR2 U333 ( .A(n622), .B(n623), .Z(n147) );
  AN2 U334 ( .A(n301), .B(n500), .Z(n623) );
  IV U335 ( .A(n302), .Z(n500) );
  AN2 U336 ( .A(n302), .B(n501), .Z(n622) );
  IV U337 ( .A(n301), .Z(n501) );
  OR2 U338 ( .A(n624), .B(n625), .Z(n119) );
  AN2 U339 ( .A(n298), .B(n520), .Z(n625) );
  IV U340 ( .A(n299), .Z(n520) );
  AN2 U341 ( .A(n299), .B(n527), .Z(n624) );
  IV U342 ( .A(n298), .Z(n527) );
  OR2 U343 ( .A(n626), .B(n627), .Z(n118) );
  AN2 U344 ( .A(n296), .B(n528), .Z(n627) );
  IV U345 ( .A(n297), .Z(n528) );
  AN2 U346 ( .A(n297), .B(n529), .Z(n626) );
  IV U347 ( .A(n296), .Z(n529) );
  OR2 U348 ( .A(n628), .B(n629), .Z(n116) );
  AN2 U349 ( .A(n28), .B(n511), .Z(n629) );
  IV U350 ( .A(n630), .Z(n628) );
  OR2 U351 ( .A(n511), .B(n28), .Z(n630) );
  AN2 U352 ( .A(n631), .B(n632), .Z(n113) );
  IV U353 ( .A(n633), .Z(n632) );
  AN2 U354 ( .A(n511), .B(n55), .Z(n633) );
  OR2 U355 ( .A(n55), .B(n511), .Z(n631) );
  IV U356 ( .A(n300), .Z(n511) );
  OR2 U357 ( .A(n634), .B(n635), .Z(U5_DATA2_5) );
  IV U358 ( .A(n636), .Z(n635) );
  OR2 U359 ( .A(n614), .B(n[9]), .Z(n636) );
  AN2 U360 ( .A(n[9]), .B(n614), .Z(n634) );
  OR2 U361 ( .A(n637), .B(n638), .Z(U5_DATA2_4) );
  IV U362 ( .A(n639), .Z(n638) );
  OR2 U363 ( .A(n614), .B(n[8]), .Z(n639) );
  AN2 U364 ( .A(n[8]), .B(n614), .Z(n637) );
  IV U365 ( .A(n21), .Z(n614) );
  OR2 U366 ( .A(n640), .B(n184), .Z(U4_Z_0) );
  AN2 U367 ( .A(CNTL_RESETN_P0), .B(n549), .Z(n640) );
  IV U368 ( .A(n293), .Z(n549) );
endmodule

