// Benchmark "Huffman_random_8" written by ABC on Fri Nov 21 18:13:42 2014

module Huffman_random_8 ( clock, 
    in_0 , in_1 , in_2 , in_3 , in_4 , in_5 , in_6 , in_7 ,
    carestate, out  );
  input  clock;
  input  in_0 , in_1 , in_2 , in_3 , in_4 , in_5 , in_6 ,
    in_7 ;
  output carestate, out;
  reg reg_0 , reg_1 , reg_2 , reg_3 , reg_4 , reg_5 , reg_6 ,
    reg_7 , counter_0 , counter_1 , counter_2 , counter_3 ,
    counter_4 ;
  wire n50, n59, n60, n61, n62_1, n63, n64, n65, n66, n67_1, n68, n69, n70,
    n71, n72_1, n73, n79, n80, n81, n82_1, n83, n84, n85, n86, n87, n88,
    n90, n91, n22, n27, n32, n37, n42, n47, n52, n57, n62, n67, n72, n77,
    n82;
  assign n50 = ~counter_0  & ~counter_1  & ~counter_2  & ~counter_3  & ~counter_4 ;
  assign n22 = n50 ? in_0  : reg_0 ;
  assign n27 = n50 ? in_1  : reg_1 ;
  assign n32 = n50 ? in_2  : reg_2 ;
  assign n37 = n50 ? in_3  : reg_3 ;
  assign n42 = n50 ? in_4  : reg_4 ;
  assign n47 = n50 ? in_5  : reg_5 ;
  assign n52 = n50 ? in_6  : reg_6 ;
  assign n57 = n50 ? in_7  : reg_7 ;
  assign n59 = in_0  & in_1  & in_2  & ~in_3  & in_4  & (in_6  ? (in_5  ^ in_7 ) : in_5 );
  assign n60 = ((in_1  ^ in_3 ) & ((~in_2  & (in_0  ? (~in_5  & (~in_4  ^ in_6 )) : (in_4  & in_5 ))) | (~in_0  & in_2  & in_4 ) | ((in_2  ? (in_6  & in_7 ) : (~in_6  & ~in_7 )) & (in_0  ? (in_4  & in_5 ) : (~in_4  & ~in_5 ))) | (~in_4  & ((~in_0  & ((in_6  & in_7  & ~in_2  & ~in_5 ) | (~in_6  & ~in_7  & in_2  & in_5 ))) | (in_0  & ~in_2  & in_5  & ~in_6  & ~in_7 ))))) | (in_0  & ((in_1  & in_3  & ~in_5  & (in_2  ^ in_4 )) | (~in_1  & ~in_3  & in_5  & (~in_2  ^ in_4 )) | (in_2  & ((~in_3  & (in_1  ? (in_4  ? (~in_5  & ~in_6 ) : (in_5  & in_6 )) : (~in_5  & ~in_6 ))) | (~in_1  & in_3  & in_4  & in_5  & ~in_6 ))) | (~in_1  & ~in_2  & ((in_3  & ~in_4  & in_6 ) | (~in_5  & ~in_6  & ~in_3  & in_4 ))))) | (~in_0  & (((~in_5  ^ ~in_6 ) & ((~in_1  & ~in_3  & (~in_2  ^ in_4 )) | (in_1  & ~in_2  & in_3  & in_4 ))) | (~in_2  & ((~in_3  & ((~in_1  & in_4  & ~in_5 ) | (in_5  & in_6  & in_1  & ~in_4 ))) | (in_1  & in_3  & in_6  & (~in_4  ^ in_5 )))) | (in_2  & ~in_4  & ~in_5  & (in_1  ? (in_3  & ~in_6 ) : ~in_3 )))) | (~in_2  & (((in_6  ^ in_7 ) & ((in_0  & in_1  & (in_3  ? (~in_4  & ~in_5 ) : (in_4  & in_5 ))) | (~in_0  & ~in_1  & in_3  & ~in_4  & ~in_5 ))) | (in_1  & ((in_7  & ((in_4  & ~in_5  & (in_0  ? (~in_3  & ~in_6 ) : (~in_3  ^ ~in_6 ))) | (in_0  & ~in_4  & in_5  & (in_3  ^ ~in_6 )))) | (~in_6  & ~in_7  & ((~in_0  & ~in_3  & (~in_4  ^ ~in_5 )) | (in_4  & in_5  & in_0  & in_3 ))))) | (in_0  & ~in_1  & ~in_3  & in_4  & ~in_5  & in_6  & ~in_7 ))) | (in_2  & ((~in_7  & (in_1  ? (in_0  ? ((~in_3  & in_4  & ~in_5  & in_6 ) | (in_5  & ~in_6  & in_3  & ~in_4 )) : (in_3  & (in_4  ? (in_5  & ~in_6 ) : (~in_5  & in_6 )))) : (in_4  & in_6  & (in_0  ? (~in_3  ^ in_5 ) : (~in_3  & in_5 ))))) | (in_6  & in_7  & ((in_0  & ~in_1  & (in_3  ? (in_4  & ~in_5 ) : (~in_4  & in_5 ))) | (in_3  & in_4  & ~in_5  & ~in_0  & in_1 )))));
  assign n61 = ((in_2  ^ ~in_5 ) & (in_3  ? (in_0  ? ((in_6  & in_7  & in_1  & ~in_4 ) | (~in_6  & ~in_7  & ~in_1  & in_4 )) : (in_1  & (in_4  ? (in_6  & in_7 ) : ~in_6 ))) : (((in_6  ^ in_7 ) & (in_0  ? (~in_1  & ~in_4 ) : in_1 )) | (~in_1  & ~in_4  & ~in_6  & (~in_0  | (in_0  & ~in_7 )))))) | (((~in_0  & ~in_4  & in_5  & in_7 ) | (in_0  & in_4  & ~in_5  & ~in_7 )) & ((in_2  & (in_1  ? (~in_3  & in_6 ) : in_3 )) | (in_1  & ~in_2  & ~in_6 ))) | ((in_2  ? (~in_5  & ~in_6 ) : (in_5  & in_6 )) & ((in_0  & in_1  & in_3 ) | (~in_0  & ~in_1  & ~in_3 ) | (~in_4  & (in_0  ? (in_1  & ~in_3 ) : (~in_1  & in_3 ))))) | (~in_4  & (in_5  ? (in_0  ? ((~in_6  & (in_1  ? (in_2  ^ in_3 ) : (in_2  & in_3 ))) | (~in_1  & in_6  & (~in_2  ^ in_3 ))) : ((in_3  & (in_1  ? in_6  : (~in_2  & ~in_6 ))) | (~in_3  & in_6  & ~in_1  & in_2 ))) : ((in_0  & ((in_6  & ((~in_1  & in_2  & in_3 ) | (~in_3  & (in_1  | (~in_1  & in_2 ))))) | (in_3  & ~in_6  & ~in_1  & in_2 ))) | (~in_0  & in_1  & in_2  & ~in_3  & ~in_6 )))) | (in_4  & (in_0  ? (~in_1  & ~in_2  & in_5  & (~in_3  | (in_3  & in_6 ))) : ((in_3  & ((~in_5  & (in_2  ? (in_1  ^ in_6 ) : ~in_1 )) | (in_5  & in_6  & ~in_1  & ~in_2 ))) | (~in_1  & ~in_2  & ~in_3  & in_5  & ~in_6 )))) | (in_6  & ((in_7  & ((in_2  & ((~in_5  & ((in_0  & ~in_1  & in_4 ) | (in_3  & ~in_4  & ~in_0  & in_1 ))) | (~in_3  & in_4  & in_5  & (~in_0  | (in_0  & in_1 ))))) | (in_0  & ~in_2  & ~in_3  & (in_1  ? (in_4  & in_5 ) : ~in_5 )))) | (in_2  & ~in_7  & ((~in_0  & ((in_3  & (in_1  ^ ~in_4 )) | (in_1  & ~in_3  & ~in_4  & ~in_5 ))) | (in_0  & in_1  & in_3  & ~in_4  & in_5 ))))) | (~in_6  & ((in_3  & ((in_7  & ((in_5  & (((in_1  ^ ~in_2 ) & (in_0  ^ in_4 )) | (in_0  & ~in_2  & in_4 ))) | (in_0  & ~in_1  & in_4  & ~in_5 ))) | (in_1  & ~in_2  & ~in_7  & (in_0  ? (~in_4  & ~in_5 ) : (in_4  | (~in_4  & in_5 )))))) | (in_0  & ~in_1  & ~in_2  & ~in_3  & in_4  & ~in_5  & ~in_7 )));
  assign n62_1 = ((~in_4  ^ ~in_5 ) & (((in_1  ? (~in_6  & in_7 ) : (in_6  & ~in_7 )) & (in_0  ? (in_2  & in_3 ) : (~in_2  & ~in_3 ))) | (~in_6  & ((in_3  & (in_0  ? (~in_1  & in_2 ) : (in_1  ^ ~in_2 ))) | (in_0  & in_2  & ~in_3 ))) | (~in_0  & ~in_1  & ~in_2  & in_3  & in_6 ) | (in_3  & (((in_0  ^ in_2 ) & (in_1  ? (in_6  & ~in_7 ) : (~in_6  & in_7 ))) | (in_1  & ~in_2  & (in_0  ? (~in_6  & in_7 ) : (in_6  & ~in_7 ))))) | (~in_0  & ~in_1  & in_2  & ~in_3  & ~in_6  & ~in_7 ))) | (in_0  & ~in_2  & ((in_3  & in_4  & in_5  & in_7 ) | (~in_5  & ~in_7  & ~in_3  & ~in_4 ))) | (~in_0  & in_2  & in_3  & in_4  & in_5  & in_7 ) | (in_7  & ((in_0  & ((~in_3  & ((in_1  & (in_2  ? (~in_4  ^ in_5 ) : (in_4  & in_5 ))) | (~in_4  & ~in_5  & ~in_1  & ~in_2 ))) | (~in_1  & in_2  & in_3  & (~in_4  ^ in_5 )))) | (in_3  & ~in_4  & ~in_5  & ~in_0  & in_1  & in_2 ))) | (~in_0  & ~in_7  & ((~in_1  & ((in_2  & in_3  & (~in_4  ^ in_5 )) | (in_4  & in_5  & ~in_2  & ~in_3 ))) | (in_1  & in_2  & ~in_3  & ~in_4  & ~in_5 ))) | (in_3  & (((in_0  ? (in_5  & in_6 ) : (~in_5  & ~in_6 )) & ((~in_1  & in_2  & (in_4  ^ in_7 )) | (in_1  & ~in_2  & in_4  & ~in_7 ))) | (~in_4  & (in_0  ? ((in_6  & ((in_1  & in_7  & (in_2  ^ ~in_5 )) | (~in_5  & ~in_7  & ~in_1  & in_2 ))) | (in_1  & ~in_2  & ~in_6  & ~in_7 )) : ((in_5  & in_6  & ~in_1  & in_2 ) | (~in_5  & ~in_6  & in_1  & ~in_2 ) | (in_1  & ((in_2  & (in_5  ? (in_6  & in_7 ) : (~in_6  & ~in_7 ))) | (~in_6  & in_7  & ~in_2  & in_5 )))))) | (in_1  & in_4  & ((~in_7  & ((~in_0  & in_5  & in_6 ) | (~in_5  & ~in_6  & in_0  & in_2 ))) | (~in_0  & ~in_2  & in_5  & ~in_6  & in_7 ))))) | (~in_3  & (in_5  ? (((in_4  ^ in_7 ) & ((in_0  & (in_1  ? (in_2  & in_6 ) : (~in_2  & ~in_6 ))) | (~in_0  & in_1  & in_2  & ~in_6 ))) | (in_6  & ((~in_7  & (in_0  ? (in_1  ? (~in_2  & in_4 ) : (in_2  & ~in_4 )) : (in_2  & ~in_4 ))) | (~in_0  & ~in_1  & in_7  & (in_2  | (~in_2  & ~in_4 ))))) | (~in_1  & ~in_2  & ~in_6  & (in_0  ? (~in_4  ^ in_7 ) : (in_4  & in_7 )))) : (in_7  ? (((~in_0  ^ in_6 ) & (in_1  ? (~in_2  & ~in_4 ) : in_4 )) | (~in_1  & ~in_4  & (in_0  ? (in_2  & in_6 ) : (~in_2  & ~in_6 )))) : ((in_6  & ((in_2  & (in_0  ? (in_1  | (~in_1  & ~in_4 )) : (~in_1  & ~in_4 ))) | (~in_0  & in_1  & ~in_2 ))) | (~in_0  & ~in_1  & ~in_2  & ~in_4  & ~in_6 )))));
  assign n63 = ((in_2  ? (~in_3  & ~in_7 ) : (in_3  & in_7 )) & (in_0  ? (in_6  ? ~in_5  : (in_1  ? (in_4  & ~in_5 ) : (~in_4  & in_5 ))) : (in_5  & (in_1  ? (in_4  | (~in_4  & in_6 )) : (in_4  & in_6 ))))) | (~in_0  & ((~in_4  & ((in_5  & ((in_1  & (in_2  ? (in_3  & ~in_6 ) : (~in_3  & in_6 ))) | (~in_3  & ~in_6  & ~in_1  & in_2 ))) | (in_3  & ~in_5  & (in_1  ? (in_2  & ~in_6 ) : ~in_2 )))) | (in_3  & in_4  & ((~in_1  & (in_2  ? in_5  : (~in_5  & ~in_6 ))) | (~in_5  & ~in_6  & in_1  & in_2 ))) | ((in_1  ^ in_3 ) & ((in_4  & ((~in_6  & in_7  & in_2  & ~in_5 ) | (in_6  & ~in_7  & ~in_2  & in_5 ))) | (in_2  & ~in_4  & in_6  & (~in_5  ^ in_7 )))) | (~in_6  & (in_5  ? (((in_2  ? (~in_3  & in_7 ) : (in_3  & ~in_7 )) & (~in_1  ^ ~in_4 )) | (~in_2  & ((~in_1  & ~in_7  & (in_3  ^ in_4 )) | (in_1  & ~in_3  & in_4  & in_7 ))) | (in_1  & in_2  & in_4  & in_7 )) : ((in_1  & ((~in_2  & (in_3  ? (in_4  ^ in_7 ) : (in_4  & in_7 ))) | (in_2  & ~in_3  & ~in_4  & in_7 ))) | (~in_1  & ~in_2  & ~in_3  & in_4  & ~in_7 )))) | (in_6  & ((in_1  & ((~in_7  & ((~in_5  & (in_2  ? (in_3  ^ in_4 ) : (~in_3  ^ in_4 ))) | (in_4  & in_5  & ~in_2  & in_3 ))) | (in_2  & in_3  & in_4  & in_5  & in_7 ))) | (in_4  & in_5  & in_7  & ~in_1  & ~in_2  & ~in_3 ))))) | (in_0  & ((~in_7  & (in_1  ? ((~in_4  & in_6  & in_2  & in_3 ) | (~in_2  & ~in_3  & in_4  & ~in_6 )) : ((~in_2  & in_4  & (in_3  ^ ~in_6 )) | (~in_4  & ~in_6  & in_2  & in_3 )))) | (~in_1  & in_7  & ((~in_6  & (in_2  ? (in_3  & in_4 ) : ~in_3 )) | (~in_4  & in_6  & ~in_2  & ~in_3 ))) | (~in_4  & (in_6  ? (((~in_2  ^ in_7 ) & (in_1  ^ ~in_5 )) | (~in_3  & ((~in_5  & in_7  & in_1  & ~in_2 ) | (in_5  & ~in_7  & ~in_1  & in_2 )))) : ((~in_3  & ((in_2  & (in_1  ? ~in_5  : (in_5  & in_7 ))) | (~in_5  & ~in_7  & ~in_1  & ~in_2 ))) | (in_1  & in_2  & in_3  & ~in_5  & ~in_7 )))) | (in_4  & ((in_2  & ((~in_5  & (((in_1  ^ in_6 ) & (in_3  ^ in_7 )) | (~in_1  & in_3  & ~in_6  & ~in_7 ))) | (in_1  & ~in_3  & in_5  & ~in_6  & ~in_7 ))) | (~in_1  & ~in_2  & (in_3  ? (~in_5  & ~in_6 ) : (in_5  & in_6 )))))));
  assign n64 = 1'b0;
  assign n65 = counter_4  | n64;
  assign n66 = counter_3  | n65;
  assign n67_1 = counter_2  | n66;
  assign n68 = counter_1  | n67_1;
  assign n69 = counter_0  ^ ~n68;
  assign n70 = counter_1  ^ ~n67_1;
  assign n71 = counter_2  ^ ~n66;
  assign n72_1 = counter_3  ^ ~n65;
  assign n73 = counter_4  ^ ~n64;
  assign n62 = n50 ? n59 : n69;
  assign n67 = n50 ? n60 : n70;
  assign n72 = n50 ? n61 : n71;
  assign n77 = n50 ? n62_1 : n72_1;
  assign n82 = n50 ? n63 : n73;
  assign n79 = in_0  ^ ~reg_0 ;
  assign n80 = in_1  ^ ~reg_1 ;
  assign n81 = in_2  ^ ~reg_2 ;
  assign n82_1 = in_3  ^ ~reg_3 ;
  assign n83 = in_4  ^ ~reg_4 ;
  assign n84 = in_5  ^ ~reg_5 ;
  assign n85 = in_6  ^ ~reg_6 ;
  assign n86 = in_7  ^ ~reg_7 ;
  assign n87 = n86 & n85 & n84 & n83 & n82_1 & n81 & n79 & n80;
  assign n88 = in_0  & in_1  & in_2  & in_3  & in_4  & (in_5  | (~in_5  & in_6 ));
  assign carestate = n50 ? ~n88 : n87;
  assign n90 = in_0  & (in_1  | (~in_1  & in_2 ) | (~in_1  & ~in_2  & in_3 ) | (~in_3  & in_4  & ~in_1  & ~in_2 ) | (~in_3  & ~in_4  & in_5  & ~in_1  & ~in_2 ) | (~in_4  & ~in_5  & in_6  & ~in_1  & ~in_2  & ~in_3 ) | (~in_1  & ~in_2  & ~in_3  & ~in_4  & ~in_5  & ~in_6  & in_7 ));
  assign n91 = ((reg_6  ^ reg_7 ) & ((~counter_0  & (reg_3  ? ((~counter_1  & counter_2  & ((~reg_0  & ((~counter_3  & (reg_1  ? (~reg_2  & reg_4 ) : (reg_2  & ~reg_4 ))) | (counter_3  & ~reg_1  & reg_2  & reg_4 ))) | (~counter_3  & reg_0  & ~reg_1  & reg_2  & ~reg_4 ))) | (counter_1  & ~counter_2  & ~counter_3  & ~reg_0  & ~reg_1  & reg_2  & reg_4 ) | (~counter_3  & ((reg_4  & ((reg_5  & ((counter_1  & ~counter_2  & (reg_0  ? (~reg_1  & reg_2 ) : (reg_1  & ~reg_2 ))) | (~counter_1  & counter_2  & ~reg_0  & reg_1  & reg_2 ))) | (~counter_1  & counter_2  & reg_0  & ~reg_1  & reg_2  & ~reg_5 ))) | (~counter_1  & counter_2  & reg_0  & reg_1  & reg_2  & ~reg_4  & reg_5 ))) | (~counter_1  & counter_3  & ((counter_2  & reg_0  & ~reg_1  & reg_2  & reg_4  & reg_5 ) | (~counter_2  & ~reg_0  & reg_1  & ~reg_2  & ~reg_4  & ~reg_5 )))) : ((reg_5  & ((reg_2  & ((reg_1  & ((reg_4  & (counter_1  ^ counter_3 ) & (counter_2  ^ reg_0 )) | (~counter_1  & counter_3  & ~reg_0  & ~reg_4 ))) | (~counter_1  & ~counter_2  & counter_3  & ~reg_1  & (reg_0  ^ reg_4 )))) | (~counter_1  & ~counter_2  & counter_3  & ~reg_2  & reg_4  & (~reg_0  ^ reg_1 )))) | (reg_1  & reg_2  & ~reg_5  & ((counter_1  & ~counter_2  & ~counter_3  & ~reg_0  & reg_4 ) | (~counter_1  & counter_2  & counter_3  & reg_0  & ~reg_4 )))))) | (counter_0  & ~counter_1  & ~counter_2  & ~counter_3  & reg_0  & reg_1  & reg_2  & ~reg_3  & reg_4  & reg_5 ) | (~counter_0  & ((counter_3  & ((reg_4  & ((~counter_2  & ((counter_1  & reg_2  & ((~counter_4  & ~reg_0  & ~reg_1  & reg_3 ) | (counter_4  & reg_0  & reg_1  & ~reg_3 ))) | (~counter_1  & counter_4  & ~reg_0  & reg_1  & ~reg_2  & ~reg_3 ))) | (~counter_1  & counter_2  & ~counter_4  & reg_1  & (reg_0  ? (~reg_2  & ~reg_3 ) : (reg_2  & reg_3 ))))) | (~counter_1  & ~counter_4  & reg_0  & reg_1  & reg_3  & ~reg_4  & (counter_2  ^ reg_2 )))) | (~counter_3  & reg_1  & ((~counter_2  & ((counter_1  & ~counter_4  & reg_0  & ~reg_2  & ~reg_3  & reg_4 ) | (~counter_1  & counter_4  & ~reg_0  & reg_2  & reg_3  & ~reg_4 ))) | (~counter_1  & counter_2  & ((~counter_4  & ((reg_0  & ~reg_3  & (reg_2  ^ reg_4 )) | (~reg_0  & ~reg_2  & reg_3  & ~reg_4 ))) | (counter_4  & ~reg_0  & reg_2  & reg_3  & ~reg_4 ))))) | (~counter_2  & ((~counter_3  & (counter_1  ? (reg_1  & ((counter_4  & ~reg_0  & ~reg_3  & reg_4  & reg_5 ) | (~counter_4  & reg_0  & reg_3  & ~reg_4  & ~reg_5 ))) : (counter_4  & reg_0  & ~reg_1  & reg_4  & (~reg_3  ^ reg_5 )))) | (~counter_1  & counter_3  & ~counter_4  & ~reg_0  & reg_4  & reg_5  & reg_1  & reg_3 ))) | (~counter_1  & counter_2  & ~reg_4  & ((counter_3  & ~counter_4  & reg_5  & (reg_0  ? (~reg_1  & ~reg_3 ) : (reg_1  & reg_3 ))) | (~counter_3  & counter_4  & reg_0  & reg_1  & reg_3  & ~reg_5 ))) | (~counter_2  & (counter_3  ? ((reg_4  & (((~reg_3  ^ ~reg_5 ) & ((~counter_1  & counter_4  & reg_2  & (~reg_0  ^ ~reg_1 )) | (counter_1  & ~counter_4  & reg_0  & reg_1  & ~reg_2 ))) | (~reg_0  & ((reg_1  & ((counter_1  & reg_5  & (counter_4  ? (~reg_2  & reg_3 ) : (reg_2  & ~reg_3 ))) | (~counter_1  & ~counter_4  & reg_2  & ~reg_3  & ~reg_5 ))) | (~counter_1  & ~reg_1  & ((reg_3  & (counter_4  ? (~reg_2  ^ reg_5 ) : (reg_2  & ~reg_5 ))) | (~counter_4  & ~reg_2  & ~reg_3  & ~reg_5 ))))) | (~counter_1  & reg_0  & ~reg_1  & ~reg_2  & (counter_4  ? (~reg_3  ^ reg_5 ) : (~reg_3  & reg_5 ))))) | (~counter_1  & ~reg_4  & (reg_0  ? (counter_4  ? (reg_1  & ~reg_5  & (reg_2  ^ reg_3 )) : (~reg_1  & ~reg_2  & reg_5 )) : ((~counter_4  & (~reg_2  ^ ~reg_5 ) & (~reg_1  ^ reg_3 )) | (counter_4  & ~reg_1  & reg_2  & reg_3  & reg_5 ))))) : ((~reg_5  & ((reg_3  & ((reg_1  & (reg_2  ^ reg_4 ) & (counter_1  ? (~counter_4  & ~reg_0 ) : (counter_4  & reg_0 ))) | (~counter_1  & counter_4  & ~reg_0  & ~reg_1  & ~reg_2  & reg_4 ))) | (~counter_1  & counter_4  & ~reg_1  & reg_2  & ~reg_3  & ~reg_4 ))) | (~reg_3  & reg_5  & ((~counter_1  & counter_4  & ~reg_2  & ~reg_4  & (~reg_0  ^ reg_1 )) | (counter_1  & ~counter_4  & ~reg_0  & ~reg_1  & reg_2  & reg_4 )))))) | (counter_2  & ((~counter_1  & (reg_0  ? (counter_3  ? ((reg_2  & ((~counter_4  & ((~reg_4  & reg_5  & reg_1  & ~reg_3 ) | (~reg_1  & reg_3  & reg_4  & ~reg_5 ))) | (counter_4  & ~reg_1  & ~reg_3  & reg_4  & reg_5 ))) | (~counter_4  & reg_1  & ~reg_2  & (reg_3  ? (reg_4  & reg_5 ) : (~reg_4  & ~reg_5 )))) : (reg_4  & reg_5  & ((reg_1  & (counter_4  ? (~reg_2  & reg_3 ) : (reg_2  & ~reg_3 ))) | (counter_4  & ~reg_1  & reg_2 )))) : (reg_2  ? (reg_4  & ((~reg_3  & ((counter_3  & (counter_4  ? (~reg_1  & reg_5 ) : (reg_1  & ~reg_5 ))) | (~counter_3  & counter_4  & reg_1  & ~reg_5 ))) | (~counter_3  & counter_4  & reg_3  & (reg_1  ^ reg_5 )))) : ((reg_4  & (reg_3  ? ((counter_3  & counter_4  & reg_1  & reg_5 ) | (~counter_3  & ~counter_4  & ~reg_1  & ~reg_5 )) : (counter_4  ? (~reg_1  & ~reg_5 ) : (reg_1  & reg_5 )))) | (~reg_1  & reg_3  & ~reg_4  & (counter_3  ? (counter_4  & ~reg_5 ) : (counter_4  ^ reg_5 ))))))) | (reg_1  & reg_2  & ~reg_3  & reg_4  & reg_5  & ~counter_4  & reg_0  & counter_1  & counter_3 ))))) | (counter_0  & ~counter_1  & ~counter_2  & counter_3  & ~counter_4  & reg_0  & reg_1  & reg_2  & ~reg_3  & reg_4  & reg_5 ))) | ((reg_5  ? (~reg_6  & ~reg_7 ) : (reg_6  & reg_7 )) & ((~counter_0  & (reg_1  ? (reg_4  ? (counter_1  ? (counter_2  ? ((~counter_3  & ~counter_4  & ~reg_0  & ~reg_2  & reg_3 ) | (counter_3  & counter_4  & reg_0  & reg_2  & ~reg_3 )) : ((~counter_3  & ((~counter_4  & (~reg_0  | (reg_0  & ~reg_2  & reg_3 ))) | (counter_4  & ~reg_0  & ~reg_2  & reg_3 ))) | (counter_3  & ~counter_4  & ~reg_0  & ~reg_2  & reg_3 ))) : (counter_4  ? (reg_0  ? ((~counter_2  & ~counter_3  & ~reg_2  & reg_3 ) | (counter_2  & counter_3  & reg_2  & ~reg_3 )) : (((counter_2  ^ counter_3 ) & (reg_2  ^ ~reg_3 )) | (counter_2  & ((reg_2  & (counter_3  | (~counter_3  & ~reg_3 ))) | (~counter_3  & ~reg_2  & reg_3 ))))) : ((counter_3  & ((counter_2  & ~reg_0  & reg_3 ) | (~counter_2  & reg_0  & ~reg_3 ) | (~counter_2  & ~reg_0  & ~reg_2  & reg_3 ))) | (counter_2  & ~counter_3  & ~reg_0  & reg_2  & ~reg_3 )))) : ((~counter_1  & ((reg_3  & ((counter_2  & ~counter_3  & (~counter_4  ^ ~reg_0 )) | (~counter_4  & reg_0  & ~counter_2  & counter_3 ))) | (~counter_2  & counter_3  & ~counter_4  & ~reg_0  & ~reg_3 ))) | (counter_1  & ~counter_2  & ~counter_3  & ~counter_4  & ~reg_0  & ~reg_3 ) | (~counter_1  & (counter_2  ? (reg_2  & (((~counter_4  ^ reg_0 ) & (counter_3  ^ ~reg_3 )) | (counter_3  & (counter_4  ? (~reg_0  & ~reg_3 ) : reg_0 )))) : (counter_3  & ~reg_2  & (counter_4  ? ~reg_0  : (reg_0  & ~reg_3 ))))) | (counter_1  & ~counter_2  & ~counter_3  & ~counter_4  & reg_0  & reg_2  & reg_3 ))) : ((reg_3  & (counter_1  ? (~counter_2  & reg_2  & reg_4  & (~counter_3  | (counter_3  & ~counter_4 ) | (counter_3  & counter_4  & reg_0 ))) : (counter_2  ? ((counter_3  & ~counter_4  & reg_0  & reg_4 ) | (~counter_3  & counter_4  & ~reg_0  & ~reg_4 ) | (reg_2  & ((counter_3  & ((counter_4  & reg_4 ) | (~counter_4  & ~reg_4 ) | (~reg_0  & (counter_4  ^ reg_4 )))) | (~counter_3  & counter_4  & reg_0  & ~reg_4 )))) : ((counter_4  & (counter_3  ? (reg_2  & (reg_0  ^ reg_4 )) : (~reg_2  & (reg_0  | (~reg_0  & ~reg_4 ))))) | (counter_3  & ~counter_4  & ~reg_0  & reg_2  & ~reg_4 ))))) | (~counter_1  & ~reg_3  & ((~reg_0  & ((~counter_3  & ((~counter_2  & counter_4  & (reg_2  ^ reg_4 )) | (counter_2  & ~counter_4  & ~reg_2  & ~reg_4 ))) | (counter_2  & counter_3  & reg_2  & reg_4 ))) | (counter_3  & reg_0  & ((~counter_2  & (counter_4  ? (reg_2  & ~reg_4 ) : (~reg_2  & reg_4 ))) | (counter_2  & ~counter_4  & reg_2  & ~reg_4 )))))))) | (counter_0  & ~counter_1  & ~counter_2  & ~counter_3  & ~counter_4  & reg_0  & reg_1  & reg_2  & ~reg_3  & reg_4 ))) | (~counter_0  & ((reg_3  & (counter_3  ? ((~counter_2  & (((reg_2  ^ reg_4 ) & ((~reg_1  & reg_5  & reg_6  & ~counter_1  & ~counter_4  & ~reg_0 ) | (counter_1  & counter_4  & reg_0  & reg_1  & ~reg_5  & ~reg_6 ))) | (counter_4  & ((reg_2  & ((~reg_5  & ((~reg_0  & ((counter_1  & (reg_1  ? (~reg_4  & ~reg_6 ) : (reg_4  & reg_6 ))) | (~counter_1  & reg_1  & ~reg_4  & reg_6 ))) | (~counter_1  & reg_0  & reg_1  & ~reg_6 ))) | (~counter_1  & reg_5  & reg_6  & (reg_0  ? ~reg_4  : (reg_1  & reg_4 ))))) | (~counter_1  & ~reg_2  & ((reg_0  & ((~reg_4  & (reg_1  ? (reg_5  & ~reg_6 ) : reg_6 )) | (~reg_5  & reg_6  & ~reg_1  & reg_4 ))) | (~reg_0  & ~reg_1  & ~reg_4  & reg_5  & reg_6 ))))) | (~counter_4  & ((~counter_1  & ((reg_4  & ((~reg_0  & reg_2  & (reg_1  ? (~reg_5  & ~reg_6 ) : (reg_5  & reg_6 ))) | (reg_0  & reg_1  & ~reg_2  & reg_5  & reg_6 ))) | (~reg_0  & ~reg_1  & ~reg_4  & ~reg_5  & (reg_2  ^ reg_6 )))) | (counter_1  & ~reg_0  & reg_1  & reg_2  & ~reg_4  & ~reg_5  & ~reg_6 ))))) | (~counter_1  & counter_2  & (reg_4  ? (~reg_5  & ((counter_4  & ((reg_0  & ~reg_1  & ~reg_2  & reg_6 ) | (~reg_0  & reg_1  & reg_2  & ~reg_6 ))) | (~counter_4  & reg_0  & reg_1  & reg_2  & ~reg_6 ))) : ((reg_0  & ~reg_1  & ~reg_2  & (counter_4  ? (~reg_5  & reg_6 ) : (~reg_5  ^ reg_6 ))) | (counter_4  & ~reg_0  & reg_1  & reg_2  & ~reg_6 ))))) : (counter_2  ? ((~counter_4  & (counter_1  ? ((~reg_0  & ~reg_1  & ~reg_2  & reg_4  & reg_5  & reg_6 ) | (reg_0  & reg_1  & reg_2  & ~reg_4  & ~reg_5  & ~reg_6 )) : ((reg_2  & (reg_0  ? (reg_4  & (reg_1  ? (~reg_5  & ~reg_6 ) : (reg_5  & reg_6 ))) : (reg_1  & ~reg_4  & (~reg_5  ^ reg_6 )))) | (~reg_0  & ~reg_1  & ~reg_2  & reg_4  & reg_5  & ~reg_6 )))) | (~counter_1  & counter_4  & reg_4  & ((~reg_5  & ~reg_6  & (reg_0  ? (reg_1  & reg_2 ) : ~reg_1 )) | (~reg_0  & ~reg_1  & ~reg_2  & reg_5  & reg_6 )))) : ((~reg_0  & ((~reg_2  & reg_6  & ((counter_1  & ~counter_4  & (reg_1  ? (~reg_4  & ~reg_5 ) : (reg_4  & reg_5 ))) | (~counter_1  & counter_4  & reg_1  & reg_4  & reg_5 ))) | (~counter_1  & counter_4  & reg_2  & reg_5  & ~reg_6  & (~reg_1  ^ reg_4 )))) | (counter_4  & reg_0  & ((reg_1  & ((~counter_1  & ((reg_2  & ~reg_6  & (reg_4  ^ reg_5 )) | (~reg_2  & ~reg_4  & ~reg_5  & reg_6 ))) | (counter_1  & ~reg_2  & reg_4  & ~reg_5  & reg_6 ))) | (~counter_1  & ~reg_1  & reg_2  & ~reg_4  & reg_5  & ~reg_6 ))))))) | (~reg_3  & (counter_4  ? (reg_2  ? (reg_4  ? ((~counter_1  & ((~counter_2  & ~counter_3  & ~reg_0  & reg_5  & reg_6 ) | (counter_2  & counter_3  & reg_0  & ~reg_5  & ~reg_6 ))) | (counter_1  & ~counter_2  & ~counter_3  & reg_0  & ~reg_5  & ~reg_6 ) | (~counter_1  & ((~counter_2  & ((counter_3  & ~reg_1  & ~reg_5  & ~reg_6 ) | (~counter_3  & reg_0  & reg_1  & reg_5  & reg_6 ))) | (~reg_1  & ~reg_5  & ~reg_6  & counter_2  & ~counter_3  & ~reg_0 )))) : ((~counter_1  & ((reg_6  & ((reg_5  & ((counter_2  & (counter_3  ? (reg_0  & reg_1 ) : (~reg_0  & ~reg_1 ))) | (~reg_0  & ~reg_1  & ~counter_2  & counter_3 ))) | (~counter_2  & ~counter_3  & reg_0  & reg_1  & ~reg_5 ))) | (counter_3  & ~reg_1  & ~reg_5  & ~reg_6  & (counter_2  | (~counter_2  & reg_0 ))))) | (counter_1  & ~counter_2  & counter_3  & ~reg_0  & ~reg_1  & ~reg_5  & ~reg_6 ))) : ((~counter_1  & ((reg_1  & ((reg_0  & ((~reg_4  & ~reg_6  & ((~reg_5  & (counter_2  | (~counter_2  & ~counter_3 ))) | (~counter_2  & counter_3  & reg_5 ))) | (~counter_2  & ~counter_3  & reg_4  & reg_5  & reg_6 ))) | (~counter_3  & ~reg_0  & ((~counter_2  & reg_4  & (~reg_5  ^ reg_6 )) | (reg_5  & reg_6  & counter_2  & ~reg_4 ))))) | (reg_0  & ~reg_1  & reg_5  & ((~reg_4  & (counter_2  ? (~counter_3  ^ reg_6 ) : (counter_3  & reg_6 ))) | (~counter_2  & counter_3  & reg_4  & ~reg_6 ))))) | (counter_1  & ~counter_2  & ~counter_3  & ~reg_0  & reg_5  & reg_6  & reg_1  & ~reg_4 ))) : ((reg_0  & (counter_2  ? (~reg_5  & ((~counter_1  & ((reg_4  & ((reg_2  & (counter_3  ? reg_6  : (reg_1  & ~reg_6 ))) | (~counter_3  & ~reg_1  & ~reg_2  & ~reg_6 ))) | (~counter_3  & reg_1  & ~reg_2  & ~reg_4  & ~reg_6 ))) | (counter_1  & counter_3  & reg_1  & reg_2  & reg_4  & reg_6 ))) : ((reg_1  & ~reg_6  & ((counter_1  & ((~counter_3  & ~reg_2  & ~reg_4  & reg_5 ) | (counter_3  & reg_2  & reg_4  & ~reg_5 ))) | (~counter_1  & counter_3  & ~reg_2  & ~reg_4  & ~reg_5 ))) | (~counter_1  & counter_3  & ~reg_1  & reg_2  & reg_4  & reg_5  & reg_6 )))) | (~counter_1  & ~reg_0  & ((~reg_5  & ~reg_6  & ((counter_3  & ((~counter_2  & ~reg_1  & reg_2  & reg_4 ) | (counter_2  & reg_1  & ~reg_2  & ~reg_4 ))) | (counter_2  & ~counter_3  & reg_2  & ~reg_4 ))) | (counter_2  & ~counter_3  & reg_1  & ~reg_2  & ~reg_4  & reg_5  & reg_6 )))))) | (reg_1  & (((counter_4  ? (~reg_5  & ~reg_7 ) : (reg_5  & reg_7 )) & ((counter_2  & ((reg_6  & ((reg_0  & reg_2  & ((~reg_3  & reg_4  & (counter_1  | (~counter_1  & ~counter_3 ))) | (~counter_1  & counter_3  & reg_3  & ~reg_4 ))) | (~counter_1  & counter_3  & ~reg_0  & ~reg_2  & reg_3  & reg_4 ))) | (~counter_1  & counter_3  & ~reg_0  & ~reg_2  & ~reg_3  & ~reg_4  & ~reg_6 ))) | (~counter_1  & ~counter_2  & counter_3  & ~reg_4  & ((~reg_0  & ~reg_3  & (reg_2  ^ ~reg_6 )) | (reg_0  & ~reg_2  & reg_3  & ~reg_6 ))))) | (((~reg_4  & reg_5  & reg_6  & reg_7 ) | (reg_4  & ~reg_5  & ~reg_6  & ~reg_7 )) & ((reg_0  & (counter_1  ? ((counter_2  & ~counter_3  & ~counter_4  & ~reg_2  & reg_3 ) | (~counter_2  & counter_3  & counter_4  & reg_2  & ~reg_3 )) : (counter_2  & counter_3  & (~counter_4  ^ reg_2 ) & reg_3 ))) | (~counter_1  & ~reg_0  & ((reg_3  & ((counter_3  & (counter_2  ? (~counter_4  & reg_2 ) : (counter_4  & ~reg_2 ))) | (counter_2  & ~counter_3  & counter_4 ))) | (counter_2  & ~counter_3  & reg_2  & ~reg_3 ))))) | (reg_4  & (counter_3  ? (reg_5  ? (((~counter_4  ^ ~reg_0 ) & ((~counter_2  & ~reg_3  & ((counter_1  & reg_2  & (~reg_6  ^ reg_7 )) | (reg_6  & reg_7  & ~counter_1  & ~reg_2 ))) | (~counter_1  & counter_2  & ~reg_2  & reg_3  & reg_6  & reg_7 ))) | (~counter_1  & ((counter_2  & ((~counter_4  & ~reg_0  & reg_2  & reg_6  & reg_7 ) | (counter_4  & reg_0  & ~reg_2  & ~reg_6  & ~reg_7 ))) | (~counter_2  & ~counter_4  & ~reg_0  & reg_6  & reg_7 ) | (reg_0  & ((~reg_3  & (counter_2  ? (reg_6  & (~counter_4  ^ reg_2 ) & reg_7 ) : (counter_4  & ~reg_6  & ~reg_7 ))) | (~counter_2  & ~counter_4  & ~reg_2  & reg_3  & ~reg_6  & ~reg_7 ))) | (counter_4  & ~reg_0  & reg_3  & reg_7  & (counter_2  ? reg_2  : (~reg_2  & reg_6 ))))) | (~counter_4  & ~reg_0  & counter_1  & ~counter_2  & reg_2  & ~reg_3  & ~reg_6  & ~reg_7 )) : ((~counter_1  & (reg_2  ? ((~reg_6  & ((counter_4  & ~reg_0  & ~reg_7  & (counter_2  ^ reg_3 )) | (~counter_2  & ~counter_4  & reg_0  & reg_7 ))) | (~reg_3  & reg_6  & reg_7  & ~counter_2  & ~counter_4  & ~reg_0 )) : (counter_2  ? ((~reg_0  & ((~reg_6  & (counter_4  ? (reg_3  ^ reg_7 ) : (reg_3  & reg_7 ))) | (reg_6  & ~reg_7  & ~counter_4  & ~reg_3 ))) | (~counter_4  & reg_0  & ~reg_3  & reg_6  & reg_7 )) : ((~reg_6  & ((~reg_3  & (counter_4  ? ~reg_7  : (~reg_0  & reg_7 ))) | (~counter_4  & ~reg_0  & reg_3  & reg_7 ))) | (counter_4  & reg_0  & reg_3  & reg_6  & reg_7 ))))) | (counter_1  & ~counter_2  & counter_4  & ~reg_0  & reg_6  & ~reg_7  & ~reg_2  & reg_3 ))) : (reg_3  ? (((~reg_5  ^ reg_7 ) & ((~counter_1  & ((counter_2  & ~counter_4  & ~reg_0  & reg_2  & reg_6 ) | (~counter_2  & counter_4  & reg_0  & ~reg_2  & ~reg_6 ))) | (counter_1  & ~counter_2  & counter_4  & ~reg_0  & ~reg_2  & reg_6 ))) | (~counter_1  & ((~reg_2  & ((counter_4  & ((reg_5  & ((reg_6  & reg_7  & (counter_2  | (~counter_2  & reg_0 ))) | (~counter_2  & ~reg_0  & ~reg_6  & ~reg_7 ))) | (counter_2  & reg_0  & ~reg_5  & ~reg_6  & reg_7 ))) | (counter_2  & ~counter_4  & ~reg_5  & ~reg_7  & (~reg_0  ^ reg_6 )))) | (counter_4  & ~reg_0  & reg_2  & reg_7  & (counter_2  ? (reg_5  & reg_6 ) : (~reg_5  & ~reg_6 )))))) : (reg_0  ? (counter_2  ? (counter_4  ? ((reg_5  & ((reg_2  & (counter_1  ? (~reg_6  ^ reg_7 ) : (reg_6  & reg_7 ))) | (~reg_6  & ~reg_7  & ~counter_1  & ~reg_2 ))) | (~counter_1  & ~reg_2  & ~reg_5  & ~reg_6  & ~reg_7 )) : (reg_6  & reg_7  & (counter_1  ? (reg_2  & ~reg_5 ) : ~reg_2 ))) : ((~reg_5  & ((counter_4  & ((~counter_1  & ~reg_7  & (reg_2  ^ reg_6 )) | (reg_6  & reg_7  & counter_1  & reg_2 ))) | (counter_1  & ~counter_4  & reg_6  & (reg_2  ^ reg_7 )))) | (counter_1  & reg_5  & ~reg_6  & (counter_4  ^ reg_2 ) & ~reg_7 ))) : ((counter_1  & ~counter_2  & ~counter_4  & (reg_5  ? (reg_6  & reg_7 ) : (~reg_6  & ~reg_7 ))) | (reg_5  & reg_6  & reg_7  & ~counter_1  & counter_2  & counter_4 ) | (reg_2  & reg_6  & ((counter_1  & reg_5  & (counter_2  ^ counter_4 ) & reg_7 ) | (~counter_1  & ~counter_2  & counter_4  & ~reg_5  & ~reg_7 ))) | (~counter_1  & ~reg_2  & ~reg_6  & ~reg_7  & (counter_2  ? (~counter_4  & ~reg_5 ) : (counter_4  & reg_5 )))))))) | (~reg_4  & (reg_7  ? (counter_4  ? (((counter_3  ? (~reg_2  & reg_3 ) : (reg_2  & ~reg_3 )) & ((counter_1  & ~counter_2  & reg_0  & reg_5  & reg_6 ) | (~counter_1  & counter_2  & ~reg_0  & ~reg_5  & ~reg_6 ))) | (~counter_1  & (counter_3  ? (reg_0  & ~reg_5  & ((~reg_2  & (counter_2  ? reg_6  : (~reg_3  & ~reg_6 ))) | (~counter_2  & reg_2  & ~reg_3  & reg_6 ))) : ((reg_0  & ((reg_5  & ((reg_2  & (counter_2  ? (~reg_3  ^ reg_6 ) : (~reg_3  & ~reg_6 ))) | (~counter_2  & ~reg_2  & (~reg_3  ^ ~reg_6 )))) | (counter_2  & ~reg_2  & reg_3  & ~reg_5  & reg_6 ))) | (~counter_2  & ~reg_0  & reg_6  & (reg_2  ? (reg_3  & ~reg_5 ) : (~reg_3  ^ ~reg_5 ))))))) : ((counter_3  & ((~counter_2  & ((reg_2  & ((reg_0  & ((counter_1  & (reg_3  ? (~reg_5  & ~reg_6 ) : (reg_5  & reg_6 ))) | (~reg_5  & reg_6  & ~counter_1  & ~reg_3 ))) | (~counter_1  & ~reg_0  & reg_3  & reg_6 ))) | (~counter_1  & ~reg_2  & ((~reg_0  & reg_3  & reg_6 ) | (reg_0  & ~reg_3  & reg_5  & ~reg_6 ))))) | (~counter_1  & counter_2  & reg_0  & reg_2  & reg_3  & reg_5  & ~reg_6 ))) | (~counter_1  & counter_2  & ~counter_3  & ((reg_0  & reg_5  & ((~reg_2  & reg_3  & ~reg_6 ) | (reg_6  & (reg_2  | (~reg_2  & ~reg_3 ))))) | (~reg_0  & ~reg_2  & reg_3  & ~reg_5  & reg_6 ))))) : (((~counter_4  ^ reg_6 ) & ((~counter_1  & counter_2  & counter_3  & ((reg_0  & ~reg_2  & reg_3  & reg_5 ) | (~reg_0  & reg_2  & ~reg_3  & ~reg_5 ))) | (counter_1  & ~counter_2  & ~counter_3  & ~reg_0  & reg_2  & reg_3  & ~reg_5 ))) | (~counter_3  & (reg_3  ? ((~reg_5  & ((reg_0  & ((~reg_6  & ((reg_2  & ((~counter_1  & counter_2  & ~counter_4 ) | (counter_4  & (counter_1  | (~counter_1  & ~counter_2 ))))) | (~counter_1  & counter_2  & ~counter_4  & ~reg_2 ))) | (counter_1  & ~counter_2  & counter_4  & reg_2  & reg_6 ))) | (~counter_1  & counter_2  & counter_4  & ~reg_0  & (reg_2  ^ reg_6 )))) | (~counter_1  & ~counter_2  & counter_4  & ~reg_0  & ~reg_2  & reg_5  & reg_6 )) : ((~counter_2  & (((reg_2  ? (reg_5  & reg_6 ) : (~reg_5  & ~reg_6 )) & (counter_1  ? (~counter_4  & reg_0 ) : (counter_4  & ~reg_0 ))) | (counter_4  & ~reg_6  & ((~counter_1  & ~reg_0  & (reg_2  | (~reg_2  & reg_5 ))) | (counter_1  & reg_0  & ~reg_2  & ~reg_5 ))))) | (~counter_1  & counter_2  & ((~reg_6  & (((~reg_0  ^ reg_2 ) & ~reg_5 ) | (~counter_4  & reg_0  & reg_2  & reg_5 ))) | (counter_4  & reg_0  & ~reg_2  & reg_5  & reg_6 )))))) | (~counter_1  & counter_3  & ~reg_5  & ((~reg_0  & (counter_2  ? ((~counter_4  & (reg_2  ? reg_6  : (reg_3  & ~reg_6 ))) | (counter_4  & ~reg_2  & ~reg_3  & reg_6 )) : ((~reg_6  & ((~reg_2  & reg_3 ) | (reg_2  & ~reg_3 ) | (~counter_4  & (reg_2  ^ ~reg_3 )))) | (~counter_4  & ~reg_2  & ~reg_3  & reg_6 )))) | (~counter_4  & reg_0  & ~reg_6  & (reg_2  ? (~counter_2  ^ reg_3 ) : counter_2 ))))))))) | (~reg_1  & ((((~reg_0  & ((reg_3  & reg_4  & ((reg_5  & reg_7  & ((counter_3  & (counter_4  ? (~reg_2  & ~reg_6 ) : (reg_2  & reg_6 ))) | (~counter_3  & counter_4  & reg_2  & reg_6 ))) | (~reg_5  & ~reg_6  & ~reg_7  & ~counter_3  & ~counter_4  & reg_2 ))) | (~counter_3  & counter_4  & reg_2  & ~reg_3  & reg_6  & ~reg_7  & ~reg_4  & ~reg_5 ))) | (~counter_3  & reg_0  & reg_5  & reg_6  & reg_7  & ((counter_4  & reg_2  & reg_3  & reg_4 ) | (~counter_4  & ~reg_2  & ~reg_3  & ~reg_4 )))) & (~counter_1  ^ ~counter_2 )) | (~counter_2  & (((reg_0  ? (~reg_3  & ~reg_5 ) : (reg_3  & reg_5 )) & ((~counter_1  & counter_4  & ((~counter_3  & reg_2  & reg_4  & reg_6  & reg_7 ) | (counter_3  & ~reg_2  & ~reg_4  & ~reg_6  & ~reg_7 ))) | (counter_1  & ~counter_3  & ~counter_4  & ~reg_2  & reg_4  & ~reg_6  & ~reg_7 ))) | (reg_4  & ((((~counter_4  & reg_5  & reg_6  & reg_7 ) | (counter_4  & ~reg_5  & ~reg_6  & ~reg_7 )) & ((~counter_1  & counter_3  & reg_0  & (reg_2  ^ ~reg_3 )) | (counter_1  & ~counter_3  & ~reg_0  & reg_2  & reg_3 ))) | (reg_6  & ((~counter_3  & (((reg_3  ? (reg_5  & reg_7 ) : (~reg_5  & ~reg_7 )) & ((counter_1  & ~counter_4  & reg_0  & reg_2 ) | (~counter_1  & counter_4  & ~reg_0  & ~reg_2 ))) | (~counter_1  & counter_4  & ((~reg_3  & ((reg_5  & (reg_0  ? reg_7  : (~reg_2  & ~reg_7 ))) | (~reg_0  & reg_2  & ~reg_5  & reg_7 ))) | (~reg_0  & reg_2  & reg_3  & ~reg_5  & reg_7 ))))) | (~counter_1  & counter_3  & (reg_0  ? ((~counter_4  & ~reg_7  & ((~reg_5  & (reg_2  | (~reg_2  & ~reg_3 ))) | (~reg_2  & reg_3  & reg_5 ))) | (counter_4  & reg_2  & ~reg_3  & reg_5  & reg_7 )) : ((reg_3  & ((reg_2  & (counter_4  ? (~reg_5  ^ reg_7 ) : (~reg_5  & reg_7 ))) | (~counter_4  & ~reg_2  & ~reg_5  & ~reg_7 ))) | (counter_4  & ~reg_2  & ~reg_3  & reg_7 )))))) | (~reg_6  & ((~counter_1  & (((~reg_3  ^ reg_5 ) & ((~counter_3  & counter_4  & ~reg_0  & reg_2  & reg_7 ) | (counter_3  & ~counter_4  & reg_0  & ~reg_2  & ~reg_7 ))) | (~reg_3  & ((reg_5  & ((~counter_3  & counter_4  & reg_0  & reg_7 ) | (counter_3  & ~counter_4  & ~reg_0  & ~reg_7 ) | (counter_3  & counter_4  & reg_0  & reg_2  & ~reg_7 ))) | (~counter_3  & counter_4  & reg_0  & ~reg_2  & ~reg_5  & ~reg_7 ))) | (counter_4  & reg_3  & ((~reg_5  & ((~reg_2  & ~reg_7  & (counter_3  | (~counter_3  & reg_0 ))) | (~counter_3  & reg_0  & reg_2  & reg_7 ))) | (~counter_3  & reg_0  & reg_2  & reg_5  & ~reg_7 ))))) | (~counter_4  & reg_0  & counter_1  & counter_3  & reg_2  & reg_3  & reg_5  & reg_7 ))))) | (~counter_1  & ~reg_4  & ((counter_3  & ~counter_4  & ~reg_3  & ((reg_0  & ~reg_2  & reg_6  & reg_7 ) | (~reg_0  & reg_2  & ~reg_6  & ~reg_7 ))) | (~counter_3  & counter_4  & ~reg_0  & ~reg_6  & reg_7  & ~reg_2  & reg_3 ) | ((~reg_3  ^ reg_7 ) & ((~counter_3  & counter_4  & reg_0  & (reg_2  ? (reg_5  & reg_6 ) : (~reg_5  & ~reg_6 ))) | (counter_3  & ~counter_4  & ~reg_0  & ~reg_2  & reg_5  & ~reg_6 ))) | (reg_0  & (reg_3  ? (reg_2  ? ((~reg_6  & ((counter_3  & ~counter_4  & (~reg_5  ^ reg_7 )) | (~counter_3  & counter_4  & ~reg_5  & ~reg_7 ))) | (~counter_3  & counter_4  & ~reg_5  & reg_6  & ~reg_7 )) : (reg_5  & ((counter_3  & ~counter_4  & (~reg_6  ^ reg_7 )) | (~counter_3  & counter_4  & reg_6  & reg_7 )))) : (~reg_7  & ((~reg_5  & ((counter_3  & ~counter_4  & (reg_2  ^ ~reg_6 )) | (~counter_3  & counter_4  & ~reg_2  & reg_6 ))) | (~counter_3  & counter_4  & reg_2  & reg_5  & ~reg_6 ))))) | (counter_4  & ~reg_0  & reg_7  & ((reg_6  & (((~reg_3  ^ reg_5 ) & (~counter_3  ^ reg_2 )) | (~reg_3  & (counter_3  ^ reg_2 ) & reg_5 ))) | (~counter_3  & ~reg_6  & (reg_2  ? (~reg_3  ^ ~reg_5 ) : (~reg_3  & ~reg_5 ))))))))) | (~counter_1  & counter_2  & (reg_3  ? (counter_4  ? (reg_2  ? ((((~reg_0  & (reg_5  ? (reg_6  & reg_7 ) : (~reg_6  & ~reg_7 ))) | (reg_6  & reg_7  & reg_0  & reg_5 )) & (~counter_3  ^ reg_4 )) | (~counter_3  & reg_4  & ~reg_6  & ~reg_7  & (reg_0  ^ reg_5 ))) : (((~reg_6  ^ reg_7 ) & ((~counter_3  & reg_0  & reg_4  & reg_5 ) | (~reg_4  & ~reg_5  & counter_3  & ~reg_0 ))) | (~counter_3  & ((~reg_6  & ((reg_0  & reg_7  & (reg_4  ^ reg_5 )) | (~reg_0  & ~reg_4  & ~reg_5  & ~reg_7 ))) | (~reg_0  & reg_4  & ~reg_5  & reg_6  & reg_7 ))))) : (reg_0  ? (reg_2  ? (((reg_5  ? (reg_6  & reg_7 ) : (~reg_6  & ~reg_7 )) & (~counter_3  ^ reg_4 )) | (~reg_5  & ~reg_6  & ~reg_7  & ~counter_3  & reg_4 )) : (counter_3  ? (~reg_7  & (reg_4  ? (~reg_5  & reg_6 ) : (reg_5  & ~reg_6 ))) : (reg_4  & ~reg_6  & reg_7 ))) : ((((~reg_4  & reg_5  & reg_6  & reg_7 ) | (reg_4  & ~reg_5  & ~reg_6  & ~reg_7 )) & (~counter_3  ^ reg_2 )) | (reg_2  & ~reg_4  & ((~counter_3  & (reg_5  ? (reg_6  & reg_7 ) : (~reg_6  & ~reg_7 ))) | (reg_6  & ~reg_7  & counter_3  & ~reg_5 )))))) : (reg_0  ? ((~reg_7  & (counter_3  ? ((~reg_5  & ((~reg_2  & ~reg_6  & (counter_4  | (~counter_4  & ~reg_4 ))) | (~counter_4  & reg_2  & ~reg_4  & reg_6 ))) | (counter_4  & reg_2  & reg_4  & reg_5  & ~reg_6 )) : (~reg_6  & (counter_4  ? (reg_2  ? (reg_4  & reg_5 ) : (~reg_4  & ~reg_5 )) : (~reg_2  & ~reg_4 ))))) | (reg_2  & reg_6  & reg_7  & ((counter_4  & reg_5 ) | (~counter_3  & ~counter_4  & reg_4  & ~reg_5 )))) : (((reg_4  ^ reg_7 ) & ((counter_3  & counter_4  & reg_2  & ~reg_5  & reg_6 ) | (~counter_3  & ~counter_4  & ~reg_2  & reg_5  & ~reg_6 ))) | (~counter_3  & ((reg_4  & ((reg_6  & reg_7  & (counter_4  ? (~reg_2  ^ reg_5 ) : (reg_2  & reg_5 ))) | (~counter_4  & ~reg_2  & ~reg_5  & ~reg_6  & ~reg_7 ))) | (~counter_4  & ~reg_4  & ((~reg_6  & reg_7  & reg_2  & reg_5 ) | (reg_6  & ~reg_7  & ~reg_2  & ~reg_5 ))))) | (counter_3  & ~counter_4  & ~reg_7  & ((reg_2  & (reg_4  ? (~reg_5  & reg_6 ) : (reg_5  & ~reg_6 ))) | (~reg_2  & reg_4  & ~reg_5  & ~reg_6 ))))))))))) | (~counter_3  & counter_4  & reg_0  & counter_0  & ~counter_1  & ~counter_2  & reg_1  & reg_2  & ~reg_3  & reg_4  & reg_5  & ~reg_6  & ~reg_7 );
  assign out = n50 ? n90 : n91;
  always @ (posedge clock) begin
    reg_0  <= n22;
    reg_1  <= n27;
    reg_2  <= n32;
    reg_3  <= n37;
    reg_4  <= n42;
    reg_5  <= n47;
    reg_6  <= n52;
    reg_7  <= n57;
    counter_0  <= n62;
    counter_1  <= n67;
    counter_2  <= n72;
    counter_3  <= n77;
    counter_4  <= n82;
  end
  initial begin
    reg_0  <= 1'b0;
    reg_1  <= 1'b0;
    reg_2  <= 1'b0;
    reg_3  <= 1'b0;
    reg_4  <= 1'b0;
    reg_5  <= 1'b0;
    reg_6  <= 1'b0;
    reg_7  <= 1'b0;
    counter_0  <= 1'b0;
    counter_1  <= 1'b0;
    counter_2  <= 1'b0;
    counter_3  <= 1'b0;
    counter_4  <= 1'b0;
  end
endmodule


