
module pcs_tx_dpath ( txclk, reset_tx, txd, tx_en, tx_er, adver_reg, ack, 
        txd_sel, tx_enc_ctrl_sel, tx_enc_conf_sel, link_up_loc, 
        jitter_study_pci, tx_10bdata, tx_en_d, tx_er_d, txd_eq_crs_ext, 
        pos_disp_tx_p, assertion_shengyushen );
  input [7:0] txd;
  input [12:0] adver_reg;
  input [1:0] txd_sel;
  input [3:0] tx_enc_ctrl_sel;
  input [3:0] tx_enc_conf_sel;
  input [1:0] jitter_study_pci;
  output [9:0] tx_10bdata;
  input txclk, reset_tx, tx_en, tx_er, ack, link_up_loc;
  output tx_en_d, tx_er_d, txd_eq_crs_ext, pos_disp_tx_p,
         assertion_shengyushen;
  wire   n3, n6, n13, n27, n28, n35, n48, n52, n55, n65, n66, n67, n68, n69,
         n70, n76, n77, n78, n79, n80, n85, n86, n87, n90, n91, n94, n99, n100,
         n103, n106, n109, n110, n113, n116, n123, n124, n125, n128, n133,
         n158, n159, n176, n191, n194, n195, n228, n229, n262, n295, n328,
         n367, n368, n397, n428, n461, n494, n495, n506, n515, n530, n545,
         n546, n565, n572, n577, n580, n585, n586, n587, n588, n589, n590,
         n593, n596, n601, n608, n609, n610, n613, n614, n615, n616, n619,
         n622, n627, n634, n635, n644, n649, n650, n653, n654, n657, n658,
         n659, n660, n661, n662, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n677, n678, n704, n705, n711, n712, n713, n738, n746,
         n747, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n997, n998, n1001, n1004, n1005, n1006, n1009, n1012,
         n1015, n1016, n1019, n1020, n1023, n1026, n1031, n1038, n1039, n1042,
         n1043, n1044, n1067, n1072, n1075, n1080, n1113, n1146, n1179, n1212,
         n1213, n1214, n1247, n1248, n1281, n1282, n1315, n1348, n1381, n1414,
         n1425, n1434, n1449, n1454, n1455, n1484, n1485, n1488, n1489, n1492,
         n1493, n1494, n1495, n1496, n1499, n1502, n1503, n1506, n1509, n1512,
         n1513, n1516, n1517, n1520, n1523, n1528, n1535, n1536, n1539, n1540,
         n1563, n1568, n1571, n1574, n1575, n1576, n1577, n1578, n1579, n1590,
         n1591, n1594, n1601, n1606, n1607, n1610, n1615, n1616, n1643, n1661,
         n1730, n1836, n1855, n1893, n1916, n1919, n1928, n1934, n1942, n1943,
         n1944, n1945, n1946, n1947, n1952, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1977, n1978, n1979, n1983, n1984, n1985, n1988, n1989, n1990, n1994,
         n1995, n1996, n2001, n2002, n2003, n2007, n2008, n2009, n2012, n2013,
         n2014, n2017, n2018, n2019, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2141, U51_Z_0, U51_Z_1, U51_Z_2,
         U51_Z_3, U51_Z_4, U51_Z_5, U51_Z_6, U51_Z_7, U50_Z_0, U50_Z_1,
         U50_Z_2, U50_Z_3, U50_Z_4, U50_Z_5, U50_Z_6, U50_Z_7, U50_CONTROL1,
         U50_DATA1_0, U50_DATA1_1, U50_DATA1_2, U50_DATA1_3, U50_DATA1_4,
         U50_DATA1_5, U50_DATA1_6, U50_DATA1_7, U49_Z_0, U48_Z_0,
         U47_DATA121_0, U20_Z_0, U20_Z_1, U20_Z_2, U20_Z_3, U20_Z_4, U20_Z_5,
         U20_Z_6, U20_Z_7, U20_Z_8, U20_Z_9, U6_Z_0, U5_Z_0, U5_Z_1, U5_Z_2,
         U5_Z_3, U5_Z_4, U5_Z_5, U5_Z_6, U5_Z_7, U5_Z_8, U5_Z_9, U5_DATA1_0,
         U5_DATA1_1, U5_DATA1_2, U5_DATA1_3, U5_DATA1_4, U5_DATA1_5,
         U5_DATA1_6, U5_DATA1_7, U5_DATA1_8, U5_DATA1_9, U4_Z_0, U4_Z_1,
         U4_Z_2, U4_Z_3, U4_DATA2_0, U4_DATA2_1, U4_DATA2_2, U4_DATA2_3, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2249, n2272, n2273,
         n2274, n2290, n2306, n2307, n2308, n2311, n2312, n2315, n2316, n2318,
         n2320, n2321, n2322, n2447, n2448, n2451, n2452, n2455, n2457, n2458,
         n2461, n2462, n2465, n2466, n2469, n2470, n2473, n2484, n2486, n2488,
         n2490, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166;
  wire   [2080:2079] n;

  IV I_09 ( .A(link_up_loc), .Z(n13) );
  OR2 C332 ( .A(n3452), .B(n27), .Z(n28) );
  IV I_07 ( .A(reset_tx), .Z(n35) );
  AN2 C272 ( .A(n2308), .B(n2307), .Z(n65) );
  AN2 C282 ( .A(n2306), .B(n2290), .Z(n66) );
  AN2 C292 ( .A(n2274), .B(n2273), .Z(n67) );
  AN2 C303 ( .A(n2272), .B(n2249), .Z(n68) );
  AN2 C312 ( .A(n65), .B(n66), .Z(n69) );
  AN2 C321 ( .A(n67), .B(n68), .Z(n70) );
  OR2 C54 ( .A(n2124), .B(n2123), .Z(n76) );
  OR2 C551 ( .A(n2122), .B(n2121), .Z(n77) );
  OR2 C571 ( .A(n2272), .B(n2249), .Z(n78) );
  OR2 C582 ( .A(n76), .B(n77), .Z(n79) );
  OR2 C591 ( .A(n614), .B(n78), .Z(n80) );
  OR2 C751 ( .A(n2120), .B(n2273), .Z(n85) );
  OR2 C761 ( .A(n2118), .B(n2249), .Z(n86) );
  OR2 C781 ( .A(n85), .B(n86), .Z(n87) );
  OR2 C86 ( .A(n2272), .B(n2117), .Z(n90) );
  OR2 C882 ( .A(n85), .B(n90), .Z(n91) );
  OR2 C992 ( .A(n85), .B(n78), .Z(n94) );
  OR2 C1151 ( .A(n2274), .B(n2119), .Z(n99) );
  OR2 C1182 ( .A(n99), .B(n86), .Z(n100) );
  OR2 C1281 ( .A(n99), .B(n90), .Z(n103) );
  OR2 C1391 ( .A(n99), .B(n78), .Z(n106) );
  OR2 C146 ( .A(n2274), .B(n2273), .Z(n109) );
  OR2 C149 ( .A(n109), .B(n588), .Z(n110) );
  OR2 C160 ( .A(n109), .B(n86), .Z(n113) );
  OR2 C1711 ( .A(n109), .B(n90), .Z(n116) );
  OR2 C198 ( .A(n2122), .B(n2290), .Z(n123) );
  OR2 C2011 ( .A(n76), .B(n123), .Z(n124) );
  OR2 C202 ( .A(n614), .B(n86), .Z(n125) );
  OR2 C212 ( .A(n614), .B(n90), .Z(n128) );
  OR2 C233 ( .A(n85), .B(n588), .Z(n133) );
  OR2 C364 ( .A(n2306), .B(n2121), .Z(n158) );
  OR2 C367 ( .A(n76), .B(n158), .Z(n159) );
  OR2 C453 ( .A(n99), .B(n588), .Z(n176) );
  OR2 C535 ( .A(n109), .B(n78), .Z(n191) );
  OR2 C541 ( .A(n2306), .B(n2290), .Z(n194) );
  OR2 C544 ( .A(n76), .B(n194), .Z(n195) );
  OR2 C731 ( .A(n2124), .B(n2307), .Z(n228) );
  OR2 C735 ( .A(n228), .B(n77), .Z(n229) );
  OR2 C912 ( .A(n228), .B(n123), .Z(n262) );
  OR2 C1104 ( .A(n228), .B(n158), .Z(n295) );
  OR2 C1297 ( .A(n228), .B(n194), .Z(n328) );
  OR2 C1530 ( .A(n2308), .B(n2123), .Z(n367) );
  OR2 C1534 ( .A(n367), .B(n77), .Z(n368) );
  OR2 C1691 ( .A(n367), .B(n123), .Z(n397) );
  OR2 C1872 ( .A(n367), .B(n158), .Z(n428) );
  OR2 C2065 ( .A(n367), .B(n194), .Z(n461) );
  OR2 C2268 ( .A(n2308), .B(n2307), .Z(n494) );
  OR2 C2272 ( .A(n494), .B(n77), .Z(n495) );
  OR2 C2330 ( .A(n85), .B(n649), .Z(n506) );
  OR2 C2378 ( .A(n99), .B(n649), .Z(n515) );
  OR2 C2465 ( .A(n494), .B(n123), .Z(n530) );
  OR2 C2551 ( .A(n2122), .B(n2290), .Z(n545) );
  OR2 C2554 ( .A(n494), .B(n545), .Z(n546) );
  OR2 C2673 ( .A(n494), .B(n158), .Z(n565) );
  OR2 C2711 ( .A(n614), .B(n609), .Z(n572) );
  OR2 C2736 ( .A(n634), .B(n649), .Z(n577) );
  OR2 C2749 ( .A(n634), .B(n653), .Z(n580) );
  OR2 C2770 ( .A(n2308), .B(n2307), .Z(n585) );
  OR2 C2771 ( .A(n2306), .B(n2121), .Z(n586) );
  OR2 C2772 ( .A(n2274), .B(n2119), .Z(n587) );
  OR2 C2773 ( .A(n2118), .B(n2117), .Z(n588) );
  OR2 C2774 ( .A(n585), .B(n586), .Z(n589) );
  OR2 C2775 ( .A(n587), .B(n588), .Z(n590) );
  OR2 C2788 ( .A(n587), .B(n649), .Z(n593) );
  OR2 C2801 ( .A(n587), .B(n653), .Z(n596) );
  OR2 C2828 ( .A(n608), .B(n588), .Z(n601) );
  OR2 C2868 ( .A(n2274), .B(n2273), .Z(n608) );
  OR2 C28691 ( .A(n2272), .B(n2249), .Z(n609) );
  OR2 C2871 ( .A(n608), .B(n609), .Z(n610) );
  OR2 C2879 ( .A(n2306), .B(n2290), .Z(n613) );
  OR2 C2880 ( .A(n2120), .B(n2119), .Z(n614) );
  OR2 C2882 ( .A(n585), .B(n613), .Z(n615) );
  OR2 C2883 ( .A(n614), .B(n588), .Z(n616) );
  OR2 C2896 ( .A(n614), .B(n649), .Z(n619) );
  OR2 C2909 ( .A(n614), .B(n653), .Z(n622) );
  OR2 C2936 ( .A(n634), .B(n588), .Z(n627) );
  OR2 C2976 ( .A(n2120), .B(n2273), .Z(n634) );
  OR2 C2979 ( .A(n634), .B(n609), .Z(n635) );
  OR2 C3035 ( .A(n587), .B(n609), .Z(n644) );
  OR2 C3062 ( .A(n2118), .B(n2249), .Z(n649) );
  OR2 C3064 ( .A(n608), .B(n649), .Z(n650) );
  OR2 C30771 ( .A(n2272), .B(n2117), .Z(n653) );
  OR2 C3079 ( .A(n608), .B(n653), .Z(n654) );
  AN2 C3082 ( .A(n2124), .B(n2123), .Z(n657) );
  AN2 C3083 ( .A(n2122), .B(n2121), .Z(n658) );
  AN2 C3084 ( .A(n2120), .B(n2119), .Z(n659) );
  AN2 C3085 ( .A(n2118), .B(n2117), .Z(n660) );
  AN2 C3086 ( .A(n657), .B(n658), .Z(n661) );
  AN2 C3087 ( .A(n659), .B(n660), .Z(n662) );
  OR2 C3636 ( .A(n677), .B(n672), .Z(n678) );
  OR2 C3670 ( .A(n704), .B(n705), .Z(n711) );
  OR2 C3672 ( .A(n712), .B(n711), .Z(n713) );
  OR2 C3697 ( .A(n3442), .B(n3441), .Z(n738) );
  AN2 C3716 ( .A(n2322), .B(n2321), .Z(n52) );
  AN2 C3720 ( .A(n2115), .B(n2320), .Z(n55) );
  AN2 C4250 ( .A(n746), .B(n2315), .Z(n665) );
  AN2 C4251 ( .A(n52), .B(n2320), .Z(n746) );
  AN2 C4252 ( .A(n52), .B(n2113), .Z(n666) );
  AN2 C4253 ( .A(n2321), .B(n2114), .Z(n667) );
  AN2 C4254 ( .A(n55), .B(n2315), .Z(n668) );
  AN2 C4255 ( .A(n55), .B(n2113), .Z(n669) );
  AN2 C4256 ( .A(n747), .B(n2315), .Z(n670) );
  AN2 C4257 ( .A(n2115), .B(n2114), .Z(n747) );
  AN2 C4258 ( .A(n2114), .B(n2113), .Z(n671) );
  AN2 C4259 ( .A(n2116), .B(n2315), .Z(n672) );
  AN2 C4260 ( .A(n2116), .B(n2113), .Z(n673) );
  AN2 C171 ( .A(n2308), .B(n2307), .Z(n983) );
  AN2 C182 ( .A(n2306), .B(n2290), .Z(n984) );
  AN2 C191 ( .A(n2274), .B(n2273), .Z(n985) );
  AN2 C201 ( .A(n2272), .B(n2249), .Z(n986) );
  AN2 C21 ( .A(n983), .B(n984), .Z(n987) );
  AN2 C22 ( .A(n985), .B(n986), .Z(n988) );
  OR2 C251 ( .A(n2124), .B(n2123), .Z(n989) );
  OR2 C26 ( .A(n2122), .B(n2121), .Z(n990) );
  OR2 C271 ( .A(n2120), .B(n2119), .Z(n991) );
  OR2 C281 ( .A(n2118), .B(n2249), .Z(n992) );
  OR2 C291 ( .A(n989), .B(n990), .Z(n993) );
  OR2 C30 ( .A(n991), .B(n992), .Z(n994) );
  OR2 C37 ( .A(n2272), .B(n2117), .Z(n997) );
  OR2 C391 ( .A(n991), .B(n997), .Z(n998) );
  OR2 C491 ( .A(n991), .B(n1015), .Z(n1001) );
  OR2 C55 ( .A(n2120), .B(n2273), .Z(n1004) );
  OR2 C561 ( .A(n2118), .B(n2117), .Z(n1005) );
  OR2 C581 ( .A(n1004), .B(n1005), .Z(n1006) );
  OR2 C68 ( .A(n1004), .B(n992), .Z(n1009) );
  OR2 C78 ( .A(n1004), .B(n997), .Z(n1012) );
  OR2 C87 ( .A(n2272), .B(n2249), .Z(n1015) );
  OR2 C891 ( .A(n1004), .B(n1015), .Z(n1016) );
  OR2 C951 ( .A(n2274), .B(n2119), .Z(n1019) );
  OR2 C98 ( .A(n1019), .B(n1005), .Z(n1020) );
  OR2 C108 ( .A(n1019), .B(n992), .Z(n1023) );
  OR2 C1181 ( .A(n1019), .B(n997), .Z(n1026) );
  OR2 C139 ( .A(n1038), .B(n1005), .Z(n1031) );
  OR2 C170 ( .A(n2274), .B(n2273), .Z(n1038) );
  OR2 C173 ( .A(n1038), .B(n1015), .Z(n1039) );
  OR2 C178 ( .A(n2122), .B(n2290), .Z(n1042) );
  OR2 C1811 ( .A(n989), .B(n1042), .Z(n1043) );
  OR2 C1821 ( .A(n991), .B(n1005), .Z(n1044) );
  OR2 C301 ( .A(n1019), .B(n1015), .Z(n1067) );
  OR2 C324 ( .A(n1038), .B(n992), .Z(n1072) );
  OR2 C336 ( .A(n1038), .B(n997), .Z(n1075) );
  OR2 C357 ( .A(n989), .B(n1213), .Z(n1080) );
  OR2 C534 ( .A(n989), .B(n1247), .Z(n1113) );
  OR2 C725 ( .A(n1212), .B(n990), .Z(n1146) );
  OR2 C902 ( .A(n1212), .B(n1042), .Z(n1179) );
  OR2 C1090 ( .A(n2124), .B(n2307), .Z(n1212) );
  OR2 C1091 ( .A(n2306), .B(n2121), .Z(n1213) );
  OR2 C1094 ( .A(n1212), .B(n1213), .Z(n1214) );
  OR2 C1284 ( .A(n2306), .B(n2290), .Z(n1247) );
  OR2 C1287 ( .A(n1212), .B(n1247), .Z(n1248) );
  OR2 C1489 ( .A(n2308), .B(n2123), .Z(n1281) );
  OR2 C1493 ( .A(n1281), .B(n990), .Z(n1282) );
  OR2 C1670 ( .A(n1281), .B(n1042), .Z(n1315) );
  OR2 C1862 ( .A(n1281), .B(n1213), .Z(n1348) );
  OR2 C2055 ( .A(n1281), .B(n1247), .Z(n1381) );
  OR2 C2262 ( .A(n1484), .B(n990), .Z(n1414) );
  OR2 C2320 ( .A(n1004), .B(n1488), .Z(n1425) );
  OR2 C2368 ( .A(n1019), .B(n1488), .Z(n1434) );
  OR2 C2455 ( .A(n1484), .B(n1042), .Z(n1449) );
  OR2 C2476 ( .A(n2122), .B(n2290), .Z(n1454) );
  OR2 C2479 ( .A(n1484), .B(n1454), .Z(n1455) );
  OR2 C2659 ( .A(n2308), .B(n2307), .Z(n1484) );
  OR2 C2663 ( .A(n1484), .B(n1213), .Z(n1485) );
  OR2 C2674 ( .A(n2118), .B(n2249), .Z(n1488) );
  OR2 C2676 ( .A(n991), .B(n1488), .Z(n1489) );
  OR2 C2683 ( .A(n2308), .B(n2307), .Z(n1492) );
  OR2 C2684 ( .A(n2306), .B(n2121), .Z(n1493) );
  OR2 C2686 ( .A(n2272), .B(n2117), .Z(n1494) );
  OR2 C2687 ( .A(n1492), .B(n1493), .Z(n1495) );
  OR2 C2688 ( .A(n991), .B(n1494), .Z(n1496) );
  OR2 C2701 ( .A(n991), .B(n1512), .Z(n1499) );
  OR2 C2710 ( .A(n2120), .B(n2273), .Z(n1502) );
  OR2 C2713 ( .A(n1502), .B(n1005), .Z(n1503) );
  OR2 C2726 ( .A(n1502), .B(n1488), .Z(n1506) );
  OR2 C2739 ( .A(n1502), .B(n1494), .Z(n1509) );
  OR2 C2751 ( .A(n2272), .B(n2249), .Z(n1512) );
  OR2 C2753 ( .A(n1502), .B(n1512), .Z(n1513) );
  OR2 C2762 ( .A(n2274), .B(n2119), .Z(n1516) );
  OR2 C2765 ( .A(n1516), .B(n1005), .Z(n1517) );
  OR2 C2778 ( .A(n1516), .B(n1488), .Z(n1520) );
  OR2 C2791 ( .A(n1516), .B(n1494), .Z(n1523) );
  OR2 C2818 ( .A(n1535), .B(n1005), .Z(n1528) );
  OR2 C2858 ( .A(n2274), .B(n2273), .Z(n1535) );
  OR2 C2861 ( .A(n1535), .B(n1512), .Z(n1536) );
  OR2 C2869 ( .A(n2306), .B(n2290), .Z(n1539) );
  OR2 C2872 ( .A(n1492), .B(n1539), .Z(n1540) );
  OR2 C3025 ( .A(n1516), .B(n1512), .Z(n1563) );
  OR2 C3054 ( .A(n1535), .B(n1488), .Z(n1568) );
  OR2 C3069 ( .A(n1535), .B(n1494), .Z(n1571) );
  AN2 C3072 ( .A(n2124), .B(n2123), .Z(n1574) );
  AN2 C3073 ( .A(n2122), .B(n2121), .Z(n1575) );
  AN2 C3074 ( .A(n2120), .B(n2119), .Z(n1576) );
  AN2 C3075 ( .A(n2118), .B(n2117), .Z(n1577) );
  AN2 C3076 ( .A(n1574), .B(n1575), .Z(n1578) );
  AN2 C3077 ( .A(n1576), .B(n1577), .Z(n1579) );
  AN2 C5522 ( .A(n2322), .B(n2321), .Z(n1590) );
  AN2 C5523 ( .A(n2320), .B(n2315), .Z(n1591) );
  OR2 C5531 ( .A(n2116), .B(n2115), .Z(n1594) );
  OR2 C5549 ( .A(n2320), .B(n2113), .Z(n1601) );
  OR2 C5555 ( .A(n2116), .B(n2321), .Z(n1606) );
  OR2 C5556 ( .A(n2320), .B(n2315), .Z(n1607) );
  OR2 C5561 ( .A(n2114), .B(n2113), .Z(n1610) );
  OR2 C5566 ( .A(n2322), .B(n2115), .Z(n1615) );
  OR2 C5567 ( .A(n2114), .B(n2315), .Z(n1616) );
  OR2 C5721 ( .A(n3448), .B(n3444), .Z(n1643) );
  OR2 C5739 ( .A(n3449), .B(n3445), .Z(n1661) );
  OR2 C5885 ( .A(n3446), .B(n3443), .Z(n1730) );
  OR2 C6002 ( .A(n3447), .B(n3443), .Z(n1836) );
  OR2 C6022 ( .A(n3447), .B(n3446), .Z(n1855) );
  OR2 C6061 ( .A(n3451), .B(n3450), .Z(n1893) );
  OR2 C6086 ( .A(n2312), .B(n2311), .Z(n1916) );
  OR2 C6090 ( .A(n2318), .B(n2316), .Z(n1919) );
  IV I_04 ( .A(reset_tx), .Z(n1928) );
  IV I_03 ( .A(reset_tx), .Z(n1934) );
  IV I_02 ( .A(txd_sel[1]), .Z(n1942) );
  IV I_110 ( .A(txd_sel[0]), .Z(n1943) );
  IV I_210 ( .A(n1944), .Z(n1945) );
  IV I_310 ( .A(n1946), .Z(n1947) );
  IV I_01 ( .A(reset_tx), .Z(n1952) );
  OR2 C128 ( .A(n2054), .B(n2049), .Z(n1965) );
  OR2 C127 ( .A(n1965), .B(n2043), .Z(n1964) );
  OR2 C126 ( .A(n1964), .B(n2038), .Z(n1963) );
  OR2 C125 ( .A(n1963), .B(n2032), .Z(n1962) );
  OR2 C124 ( .A(n1962), .B(n2025), .Z(n1961) );
  AN2 C123 ( .A(n2062), .B(n2060), .Z(n1968) );
  AN2 C122 ( .A(n1968), .B(link_up_loc), .Z(n1967) );
  AN2 C121 ( .A(n1967), .B(n2058), .Z(n1966) );
  AN2 C120 ( .A(n1966), .B(n1961), .Z(assertion_shengyushen) );
  AN2 C119 ( .A(tx_er_d), .B(n2215), .Z(txd_eq_crs_ext) );
  OR2 C118 ( .A(n2205), .B(n2206), .Z(n1975) );
  OR2 C117 ( .A(n1975), .B(n2207), .Z(n1974) );
  OR2 C116 ( .A(n1974), .B(n2208), .Z(n1973) );
  OR2 C115 ( .A(n1973), .B(n2209), .Z(n1972) );
  OR2 C114 ( .A(n1972), .B(n2210), .Z(n1971) );
  OR2 C113 ( .A(n1971), .B(n2211), .Z(n1970) );
  OR2 C112 ( .A(n1970), .B(n2202), .Z(n1969) );
  OR2 C111 ( .A(n1969), .B(n2203), .Z(n2141) );
  OR2 C107 ( .A(n2214), .B(n1978), .Z(n1977) );
  OR2 C106 ( .A(U4_Z_1), .B(n1979), .Z(n1978) );
  OR2 C105 ( .A(U4_Z_2), .B(n2204), .Z(n1979) );
  OR2 C101 ( .A(U4_Z_0), .B(n1984), .Z(n1983) );
  OR2 C100 ( .A(U4_Z_1), .B(n1985), .Z(n1984) );
  OR2 C99 ( .A(U4_Z_2), .B(n2204), .Z(n1985) );
  OR2 C96 ( .A(U4_Z_0), .B(n1989), .Z(n1988) );
  OR2 C95 ( .A(n2213), .B(n1990), .Z(n1989) );
  OR2 C94 ( .A(n2212), .B(U4_Z_3), .Z(n1990) );
  OR2 C90 ( .A(n2214), .B(n1995), .Z(n1994) );
  OR2 C89 ( .A(n2213), .B(n1996), .Z(n1995) );
  OR2 C88 ( .A(n2212), .B(U4_Z_3), .Z(n1996) );
  OR2 C83 ( .A(n2214), .B(n2002), .Z(n2001) );
  OR2 C82 ( .A(U4_Z_1), .B(n2003), .Z(n2002) );
  OR2 C81 ( .A(n2212), .B(U4_Z_3), .Z(n2003) );
  OR2 C77 ( .A(U4_Z_0), .B(n2008), .Z(n2007) );
  OR2 C76 ( .A(U4_Z_1), .B(n2009), .Z(n2008) );
  OR2 C75 ( .A(n2212), .B(U4_Z_3), .Z(n2009) );
  OR2 C72 ( .A(U4_Z_0), .B(n2013), .Z(n2012) );
  OR2 C71 ( .A(n2213), .B(n2014), .Z(n2013) );
  OR2 C70 ( .A(U4_Z_2), .B(U4_Z_3), .Z(n2014) );
  OR2 C67 ( .A(n2214), .B(n2018), .Z(n2017) );
  OR2 C66 ( .A(U4_Z_1), .B(n2019), .Z(n2018) );
  OR2 C65 ( .A(U4_Z_2), .B(U4_Z_3), .Z(n2019) );
  OR2 C62 ( .A(U4_Z_0), .B(n2023), .Z(n2022) );
  OR2 C61 ( .A(U4_Z_1), .B(n2024), .Z(n2023) );
  OR2 C60 ( .A(U4_Z_2), .B(U4_Z_3), .Z(n2024) );
  IV I_22 ( .A(n2026), .Z(n2025) );
  OR2 C58 ( .A(n2029), .B(n2027), .Z(n2026) );
  OR2 C57 ( .A(n2030), .B(n2028), .Z(n2027) );
  OR2 C56 ( .A(n2031), .B(tx_enc_ctrl_sel[3]), .Z(n2028) );
  IV I_21 ( .A(tx_enc_ctrl_sel[0]), .Z(n2029) );
  IV I_20 ( .A(tx_enc_ctrl_sel[1]), .Z(n2030) );
  IV I_19 ( .A(tx_enc_ctrl_sel[2]), .Z(n2031) );
  IV I_18 ( .A(n2033), .Z(n2032) );
  OR2 C51 ( .A(n2036), .B(n2034), .Z(n2033) );
  OR2 C50 ( .A(tx_enc_ctrl_sel[1]), .B(n2035), .Z(n2034) );
  OR2 C49 ( .A(n2037), .B(tx_enc_ctrl_sel[3]), .Z(n2035) );
  IV I_17 ( .A(tx_enc_ctrl_sel[0]), .Z(n2036) );
  IV I_16 ( .A(tx_enc_ctrl_sel[2]), .Z(n2037) );
  IV I_15 ( .A(n2039), .Z(n2038) );
  OR2 C45 ( .A(tx_enc_ctrl_sel[0]), .B(n2040), .Z(n2039) );
  OR2 C44 ( .A(tx_enc_ctrl_sel[1]), .B(n2041), .Z(n2040) );
  OR2 C43 ( .A(n2042), .B(tx_enc_ctrl_sel[3]), .Z(n2041) );
  IV I_14 ( .A(tx_enc_ctrl_sel[2]), .Z(n2042) );
  IV I_13 ( .A(n2044), .Z(n2043) );
  OR2 C40 ( .A(n2047), .B(n2045), .Z(n2044) );
  OR2 C39 ( .A(n2048), .B(n2046), .Z(n2045) );
  OR2 C38 ( .A(tx_enc_ctrl_sel[2]), .B(tx_enc_ctrl_sel[3]), .Z(n2046) );
  IV I_12 ( .A(tx_enc_ctrl_sel[0]), .Z(n2047) );
  IV I_11 ( .A(tx_enc_ctrl_sel[1]), .Z(n2048) );
  IV I_10 ( .A(n2050), .Z(n2049) );
  OR2 C34 ( .A(tx_enc_ctrl_sel[0]), .B(n2051), .Z(n2050) );
  OR2 C33 ( .A(n2053), .B(n2052), .Z(n2051) );
  OR2 C32 ( .A(tx_enc_ctrl_sel[2]), .B(tx_enc_ctrl_sel[3]), .Z(n2052) );
  IV I_9 ( .A(tx_enc_ctrl_sel[1]), .Z(n2053) );
  IV I_8 ( .A(n2055), .Z(n2054) );
  OR2 C29 ( .A(tx_enc_ctrl_sel[0]), .B(n2056), .Z(n2055) );
  OR2 C28 ( .A(tx_enc_ctrl_sel[1]), .B(n2057), .Z(n2056) );
  OR2 C27 ( .A(tx_enc_ctrl_sel[2]), .B(tx_enc_ctrl_sel[3]), .Z(n2057) );
  IV I_7 ( .A(n2059), .Z(n2058) );
  OR2 C25 ( .A(jitter_study_pci[0]), .B(jitter_study_pci[1]), .Z(n2059) );
  IV I_6 ( .A(n2061), .Z(n2060) );
  OR2 C23 ( .A(txd_sel[0]), .B(txd_sel[1]), .Z(n2061) );
  IV I_5 ( .A(reset_tx), .Z(n2062) );
  OR2 C20 ( .A(n2216), .B(n2065), .Z(n2064) );
  OR2 C19 ( .A(n2217), .B(n2066), .Z(n2065) );
  OR2 C18 ( .A(n2218), .B(n2067), .Z(n2066) );
  OR2 C17 ( .A(n2219), .B(n2068), .Z(n2067) );
  OR2 C16 ( .A(U50_DATA1_4), .B(n2069), .Z(n2068) );
  OR2 C15 ( .A(U50_DATA1_5), .B(n2070), .Z(n2069) );
  OR2 C14 ( .A(U50_DATA1_6), .B(U50_DATA1_7), .Z(n2070) );
  FD1 qout_reg_0_ ( .D(U51_Z_0), .CP(txclk), .Q(U50_DATA1_0) );
  FD1 qout_reg_1_ ( .D(U51_Z_1), .CP(txclk), .Q(U50_DATA1_1) );
  FD1 qout_reg_2_ ( .D(U51_Z_2), .CP(txclk), .Q(U50_DATA1_2) );
  FD1 qout_reg_3_ ( .D(U51_Z_3), .CP(txclk), .Q(U50_DATA1_3) );
  FD1 qout_reg_4_ ( .D(U51_Z_4), .CP(txclk), .Q(U50_DATA1_4) );
  FD1 qout_reg_5_ ( .D(U51_Z_5), .CP(txclk), .Q(U50_DATA1_5) );
  FD1 qout_reg_6_ ( .D(U51_Z_6), .CP(txclk), .Q(U50_DATA1_6) );
  FD1 qout_reg_7_ ( .D(U51_Z_7), .CP(txclk), .Q(U50_DATA1_7) );
  FD1 qout_reg_0_1 ( .D(U50_Z_0), .CP(txclk), .Q(n2117) );
  FD1 qout_reg_1_1 ( .D(U50_Z_1), .CP(txclk), .Q(n2118) );
  FD1 qout_reg_2_1 ( .D(U50_Z_2), .CP(txclk), .Q(n2119) );
  FD1 qout_reg_3_1 ( .D(U50_Z_3), .CP(txclk), .Q(n2120) );
  FD1 qout_reg_4_1 ( .D(U50_Z_4), .CP(txclk), .Q(n2121) );
  FD1 qout_reg_5_1 ( .D(U50_Z_5), .CP(txclk), .Q(n2122) );
  FD1 qout_reg_6_1 ( .D(U50_Z_6), .CP(txclk), .Q(n2123) );
  FD1 qout_reg_7_1 ( .D(U50_Z_7), .CP(txclk), .Q(n2124) );
  FD1 qout_reg_0_2 ( .D(U49_Z_0), .CP(txclk), .Q(tx_en_d) );
  FD1 qout_reg_0_3 ( .D(U48_Z_0), .CP(txclk), .Q(tx_er_d) );
  FD1 qout_reg_0_4 ( .D(reset_tx), .CP(txclk), .Q(n48) );
  FD1 qout_reg_0_8 ( .D(tx_enc_ctrl_sel[0]), .CP(txclk), .Q(U4_DATA2_0) );
  FD1 qout_reg_1_4 ( .D(tx_enc_ctrl_sel[1]), .CP(txclk), .Q(U4_DATA2_1) );
  FD1 qout_reg_2_4 ( .D(tx_enc_ctrl_sel[2]), .CP(txclk), .Q(U4_DATA2_2) );
  FD1 qout_reg_3_4 ( .D(tx_enc_ctrl_sel[3]), .CP(txclk), .Q(U4_DATA2_3) );
  FD1 qout_reg_0_9 ( .D(U4_Z_0), .CP(txclk), .Q(n2113) );
  FD1 qout_reg_1_5 ( .D(U4_Z_1), .CP(txclk), .Q(n2114) );
  FD1 qout_reg_2_5 ( .D(U4_Z_2), .CP(txclk), .Q(n2115) );
  FD1 qout_reg_3_5 ( .D(U4_Z_3), .CP(txclk), .Q(n2116) );
  FD1 qout_reg_0_10 ( .D(n2141), .CP(txclk), .Q(n2112) );
  FD1 qout_reg_0_5 ( .D(U6_Z_0), .CP(txclk), .Q(U47_DATA121_0) );
  FD1 qout_reg_0_6 ( .D(U20_Z_0), .CP(txclk), .Q(U5_DATA1_0) );
  FD1 qout_reg_1_2 ( .D(U20_Z_1), .CP(txclk), .Q(U5_DATA1_1) );
  FD1 qout_reg_2_2 ( .D(U20_Z_2), .CP(txclk), .Q(U5_DATA1_2) );
  FD1 qout_reg_3_2 ( .D(U20_Z_3), .CP(txclk), .Q(U5_DATA1_3) );
  FD1 qout_reg_4_2 ( .D(U20_Z_4), .CP(txclk), .Q(U5_DATA1_4) );
  FD1 qout_reg_5_2 ( .D(U20_Z_5), .CP(txclk), .Q(U5_DATA1_5) );
  FD1 qout_reg_6_2 ( .D(U20_Z_6), .CP(txclk), .Q(U5_DATA1_6) );
  FD1 qout_reg_7_2 ( .D(U20_Z_7), .CP(txclk), .Q(U5_DATA1_7) );
  FD1 qout_reg_8_ ( .D(U20_Z_8), .CP(txclk), .Q(U5_DATA1_8) );
  FD1 qout_reg_9_ ( .D(U20_Z_9), .CP(txclk), .Q(U5_DATA1_9) );
  FD1 sync1_reg ( .D(jitter_study_pci[1]), .CP(txclk), .Q(n6) );
  FD1 Q_reg ( .D(n6), .CP(txclk), .Q(n[2080]) );
  FD1 sync1_reg1 ( .D(jitter_study_pci[0]), .CP(txclk), .Q(n3) );
  FD1 Q_reg1 ( .D(n3), .CP(txclk), .Q(n[2079]) );
  FD1 qout_reg_9_1 ( .D(U5_Z_9), .CP(txclk), .Q(tx_10bdata[9]) );
  FD1 qout_reg_8_1 ( .D(U5_Z_8), .CP(txclk), .Q(tx_10bdata[8]) );
  FD1 qout_reg_2_3 ( .D(U5_Z_2), .CP(txclk), .Q(tx_10bdata[2]) );
  FD1 qout_reg_1_3 ( .D(U5_Z_1), .CP(txclk), .Q(tx_10bdata[1]) );
  FD1 qout_reg_0_7 ( .D(U5_Z_0), .CP(txclk), .Q(tx_10bdata[0]) );
  FD1 qout_reg_7_3 ( .D(U5_Z_7), .CP(txclk), .Q(tx_10bdata[7]) );
  FD1 qout_reg_5_3 ( .D(U5_Z_5), .CP(txclk), .Q(tx_10bdata[5]) );
  FD1 qout_reg_3_3 ( .D(U5_Z_3), .CP(txclk), .Q(tx_10bdata[3]) );
  FD1 qout_reg_4_3 ( .D(U5_Z_4), .CP(txclk), .Q(tx_10bdata[4]) );
  FD1 qout_reg_6_3 ( .D(U5_Z_6), .CP(txclk), .Q(tx_10bdata[6]) );
  OR2 U169 ( .A(n1942), .B(txd_sel[0]), .Z(n1946) );
  OR2 U170 ( .A(n1943), .B(txd_sel[1]), .Z(n1944) );
  AN2 U245 ( .A(n1952), .B(txd[7]), .Z(U51_Z_7) );
  AN2 U246 ( .A(txd[6]), .B(n1952), .Z(U51_Z_6) );
  AN2 U247 ( .A(txd[5]), .B(n1952), .Z(U51_Z_5) );
  AN2 U248 ( .A(txd[4]), .B(n1952), .Z(U51_Z_4) );
  AN2 U249 ( .A(txd[3]), .B(n1952), .Z(U51_Z_3) );
  AN2 U250 ( .A(txd[2]), .B(n1952), .Z(U51_Z_2) );
  AN2 U251 ( .A(txd[1]), .B(n1952), .Z(U51_Z_1) );
  AN2 U252 ( .A(txd[0]), .B(n1952), .Z(U51_Z_0) );
  AN2 U254 ( .A(n1945), .B(adver_reg[7]), .Z(n2447) );
  AN2 U258 ( .A(adver_reg[6]), .B(n1945), .Z(n2451) );
  AN2 U260 ( .A(n1947), .B(ack), .Z(n2448) );
  AN2 U263 ( .A(adver_reg[5]), .B(n1945), .Z(n2455) );
  AN2 U265 ( .A(adver_reg[12]), .B(n1947), .Z(n2452) );
  AN2 U267 ( .A(adver_reg[4]), .B(n1945), .Z(n2457) );
  AN2 U271 ( .A(adver_reg[3]), .B(n1945), .Z(n2461) );
  AN2 U273 ( .A(adver_reg[11]), .B(n1947), .Z(n2458) );
  AN2 U276 ( .A(adver_reg[2]), .B(n1945), .Z(n2465) );
  AN2 U278 ( .A(adver_reg[10]), .B(n1947), .Z(n2462) );
  AN2 U281 ( .A(adver_reg[1]), .B(n1945), .Z(n2469) );
  AN2 U283 ( .A(adver_reg[9]), .B(n1947), .Z(n2466) );
  AN2 U286 ( .A(adver_reg[0]), .B(n1945), .Z(n2473) );
  AN2 U288 ( .A(adver_reg[8]), .B(n1947), .Z(n2470) );
  AN2 U290 ( .A(n1942), .B(n1943), .Z(U50_CONTROL1) );
  AN2 U311 ( .A(n1934), .B(tx_en), .Z(U49_Z_0) );
  AN2 U312 ( .A(n1928), .B(tx_er), .Z(U48_Z_0) );
  AN2 U315 ( .A(n13), .B(tx_enc_conf_sel[3]), .Z(n2484) );
  AN2 U318 ( .A(tx_enc_conf_sel[2]), .B(n13), .Z(n2486) );
  AN2 U321 ( .A(tx_enc_conf_sel[1]), .B(n13), .Z(n2488) );
  AN2 U324 ( .A(tx_enc_conf_sel[0]), .B(n13), .Z(n2490) );
  OR2 U1295 ( .A(n3453), .B(n3454), .Z(n712) );
  OR2 U1296 ( .A(n3455), .B(n3456), .Z(n3454) );
  OR2 U1297 ( .A(n3457), .B(n3458), .Z(n3456) );
  AN2 U1298 ( .A(n70), .B(n69), .Z(n3458) );
  AN2 U1299 ( .A(n3459), .B(n3460), .Z(n3457) );
  OR2 U1300 ( .A(n3461), .B(n3462), .Z(n3455) );
  OR2 U1301 ( .A(n3463), .B(n3464), .Z(n3462) );
  AN2 U1302 ( .A(n3465), .B(n3466), .Z(n3464) );
  AN2 U1303 ( .A(n3467), .B(n3468), .Z(n3463) );
  OR2 U1304 ( .A(n3469), .B(n3470), .Z(n3467) );
  OR2 U1305 ( .A(n3471), .B(n3472), .Z(n3470) );
  AN2 U1306 ( .A(n3473), .B(n3474), .Z(n3461) );
  OR2 U1307 ( .A(n3475), .B(n3476), .Z(n3453) );
  OR2 U1308 ( .A(n3477), .B(n3478), .Z(n3476) );
  IV U1309 ( .A(n3479), .Z(n3478) );
  OR2 U1310 ( .A(n3480), .B(n495), .Z(n3479) );
  AN2 U1311 ( .A(n3481), .B(n3482), .Z(n3480) );
  AN2 U1312 ( .A(n580), .B(n80), .Z(n3482) );
  AN2 U1313 ( .A(n3483), .B(n515), .Z(n3481) );
  AN2 U1314 ( .A(n506), .B(n3484), .Z(n3483) );
  IV U1315 ( .A(n3485), .Z(n3484) );
  AN2 U1316 ( .A(n3486), .B(n3487), .Z(n3477) );
  OR2 U1317 ( .A(n3488), .B(n3489), .Z(n3475) );
  OR2 U1318 ( .A(n3490), .B(n3491), .Z(n3489) );
  AN2 U1319 ( .A(n3492), .B(n3493), .Z(n3491) );
  OR2 U1320 ( .A(n3494), .B(n3495), .Z(n3492) );
  AN2 U1321 ( .A(n3496), .B(n3497), .Z(n3490) );
  OR2 U1322 ( .A(n3498), .B(n3499), .Z(n3496) );
  AN2 U1323 ( .A(n3500), .B(n3501), .Z(n3488) );
  OR2 U1324 ( .A(n3495), .B(n3502), .Z(n3500) );
  IV U1325 ( .A(n565), .Z(n3495) );
  OR2 U1326 ( .A(n3503), .B(n3504), .Z(n705) );
  AN2 U1327 ( .A(n662), .B(n661), .Z(n3504) );
  AN2 U1328 ( .A(n3505), .B(n3506), .Z(n3503) );
  OR2 U1329 ( .A(n3507), .B(n3508), .Z(n704) );
  AN2 U1330 ( .A(n3509), .B(n3506), .Z(n3508) );
  OR2 U1331 ( .A(n3510), .B(n3493), .Z(n3509) );
  AN2 U1332 ( .A(n3511), .B(n3487), .Z(n3507) );
  OR2 U1333 ( .A(n3512), .B(n3513), .Z(n3511) );
  OR2 U1334 ( .A(n3514), .B(n3515), .Z(n677) );
  OR2 U1335 ( .A(n668), .B(n667), .Z(n3515) );
  OR2 U1336 ( .A(n669), .B(n3516), .Z(n3514) );
  OR2 U1337 ( .A(n671), .B(n670), .Z(n3516) );
  AN2 U1338 ( .A(n[2080]), .B(n3517), .Z(n3452) );
  AN2 U1339 ( .A(n3471), .B(n3506), .Z(n3442) );
  AN2 U1340 ( .A(n3472), .B(n3506), .Z(n3441) );
  AN2 U1341 ( .A(n[2079]), .B(n[2080]), .Z(n27) );
  IV U1342 ( .A(n2116), .Z(n2322) );
  IV U1343 ( .A(n2115), .Z(n2321) );
  IV U1344 ( .A(n2114), .Z(n2320) );
  IV U1345 ( .A(n2113), .Z(n2315) );
  IV U1346 ( .A(n2124), .Z(n2308) );
  IV U1347 ( .A(n2123), .Z(n2307) );
  IV U1348 ( .A(n2122), .Z(n2306) );
  IV U1349 ( .A(n2121), .Z(n2290) );
  IV U1350 ( .A(n2120), .Z(n2274) );
  IV U1351 ( .A(n2119), .Z(n2273) );
  IV U1352 ( .A(n2118), .Z(n2272) );
  IV U1353 ( .A(n2117), .Z(n2249) );
  IV U1354 ( .A(U50_DATA1_3), .Z(n2219) );
  IV U1355 ( .A(U50_DATA1_2), .Z(n2218) );
  IV U1356 ( .A(U50_DATA1_1), .Z(n2217) );
  IV U1357 ( .A(U50_DATA1_0), .Z(n2216) );
  IV U1358 ( .A(n2064), .Z(n2215) );
  IV U1359 ( .A(U4_Z_0), .Z(n2214) );
  IV U1360 ( .A(U4_Z_1), .Z(n2213) );
  IV U1361 ( .A(U4_Z_2), .Z(n2212) );
  IV U1362 ( .A(n1988), .Z(n2211) );
  IV U1363 ( .A(n1994), .Z(n2210) );
  IV U1364 ( .A(n2001), .Z(n2209) );
  IV U1365 ( .A(n2007), .Z(n2208) );
  IV U1366 ( .A(n2012), .Z(n2207) );
  IV U1367 ( .A(n2017), .Z(n2206) );
  IV U1368 ( .A(n2022), .Z(n2205) );
  IV U1369 ( .A(U4_Z_3), .Z(n2204) );
  IV U1370 ( .A(n1977), .Z(n2203) );
  IV U1371 ( .A(n1983), .Z(n2202) );
  AN2 U1372 ( .A(n35), .B(pos_disp_tx_p), .Z(U6_Z_0) );
  AN2 U1373 ( .A(n3518), .B(n3519), .Z(pos_disp_tx_p) );
  OR2 U1374 ( .A(n3520), .B(n3521), .Z(n3519) );
  OR2 U1375 ( .A(n3522), .B(n3523), .Z(n3521) );
  AN2 U1376 ( .A(n3524), .B(n3525), .Z(n3523) );
  OR2 U1377 ( .A(n665), .B(n3526), .Z(n3525) );
  OR2 U1378 ( .A(n673), .B(n666), .Z(n3526) );
  AN2 U1379 ( .A(n3527), .B(n3528), .Z(n3522) );
  AN2 U1380 ( .A(n3529), .B(n3530), .Z(n3527) );
  OR2 U1381 ( .A(n713), .B(n3531), .Z(n3530) );
  OR2 U1382 ( .A(U47_DATA121_0), .B(n3532), .Z(n3529) );
  OR2 U1383 ( .A(n3533), .B(n3534), .Z(n3532) );
  OR2 U1384 ( .A(n3535), .B(n3536), .Z(n3534) );
  OR2 U1385 ( .A(n3537), .B(n3538), .Z(n3536) );
  AN2 U1386 ( .A(n3502), .B(n3493), .Z(n3538) );
  IV U1387 ( .A(n530), .Z(n3502) );
  AN2 U1388 ( .A(n3539), .B(n3487), .Z(n3537) );
  IV U1389 ( .A(n589), .Z(n3487) );
  OR2 U1390 ( .A(n3485), .B(n3540), .Z(n3539) );
  OR2 U1391 ( .A(n3541), .B(n3542), .Z(n3485) );
  OR2 U1392 ( .A(n3472), .B(n3543), .Z(n3542) );
  IV U1393 ( .A(n601), .Z(n3472) );
  OR2 U1394 ( .A(n3505), .B(n3471), .Z(n3541) );
  IV U1395 ( .A(n596), .Z(n3471) );
  OR2 U1396 ( .A(n3544), .B(n3545), .Z(n3535) );
  OR2 U1397 ( .A(n3546), .B(n3547), .Z(n3545) );
  AN2 U1398 ( .A(n3497), .B(n3474), .Z(n3547) );
  IV U1399 ( .A(n3548), .Z(n3474) );
  AN2 U1400 ( .A(n3549), .B(n3550), .Z(n3548) );
  AN2 U1401 ( .A(n3551), .B(n103), .Z(n3550) );
  AN2 U1402 ( .A(n100), .B(n80), .Z(n3551) );
  AN2 U1403 ( .A(n3552), .B(n91), .Z(n3549) );
  AN2 U1404 ( .A(n87), .B(n110), .Z(n3552) );
  OR2 U1405 ( .A(n3494), .B(n3553), .Z(n3497) );
  OR2 U1406 ( .A(n3554), .B(n3555), .Z(n3494) );
  OR2 U1407 ( .A(n3556), .B(n3557), .Z(n3555) );
  AN2 U1408 ( .A(n3465), .B(n3460), .Z(n3546) );
  OR2 U1409 ( .A(n3558), .B(n3559), .Z(n3465) );
  OR2 U1410 ( .A(n3556), .B(n3554), .Z(n3559) );
  IV U1411 ( .A(n397), .Z(n3554) );
  IV U1412 ( .A(n124), .Z(n3556) );
  AN2 U1413 ( .A(n3459), .B(n3466), .Z(n3544) );
  IV U1414 ( .A(n3560), .Z(n3466) );
  AN2 U1415 ( .A(n3561), .B(n3562), .Z(n3560) );
  AN2 U1416 ( .A(n113), .B(n106), .Z(n3562) );
  AN2 U1417 ( .A(n94), .B(n116), .Z(n3561) );
  OR2 U1418 ( .A(n3563), .B(n3564), .Z(n3459) );
  OR2 U1419 ( .A(n3557), .B(n3553), .Z(n3564) );
  IV U1420 ( .A(n79), .Z(n3553) );
  IV U1421 ( .A(n368), .Z(n3557) );
  OR2 U1422 ( .A(n3565), .B(n3566), .Z(n3533) );
  OR2 U1423 ( .A(n3567), .B(n3568), .Z(n3566) );
  AN2 U1424 ( .A(n3569), .B(n3468), .Z(n3568) );
  IV U1425 ( .A(n546), .Z(n3468) );
  OR2 U1426 ( .A(n3510), .B(n3570), .Z(n3569) );
  OR2 U1427 ( .A(n3505), .B(n3513), .Z(n3570) );
  IV U1428 ( .A(n3571), .Z(n3505) );
  AN2 U1429 ( .A(n3572), .B(n654), .Z(n3571) );
  AN2 U1430 ( .A(n650), .B(n644), .Z(n3572) );
  OR2 U1431 ( .A(n3543), .B(n3512), .Z(n3510) );
  IV U1432 ( .A(n590), .Z(n3512) );
  IV U1433 ( .A(n635), .Z(n3543) );
  AN2 U1434 ( .A(n3573), .B(n3574), .Z(n3567) );
  IV U1435 ( .A(n495), .Z(n3574) );
  OR2 U1436 ( .A(n3460), .B(n3575), .Z(n3573) );
  OR2 U1437 ( .A(n3513), .B(n3576), .Z(n3575) );
  IV U1438 ( .A(n610), .Z(n3513) );
  IV U1439 ( .A(n3577), .Z(n3460) );
  AN2 U1440 ( .A(n3578), .B(n133), .Z(n3577) );
  AN2 U1441 ( .A(n128), .B(n125), .Z(n3578) );
  OR2 U1442 ( .A(n3579), .B(n3580), .Z(n3565) );
  OR2 U1443 ( .A(n738), .B(n3581), .Z(n3580) );
  AN2 U1444 ( .A(n3582), .B(n3473), .Z(n3581) );
  OR2 U1445 ( .A(n3558), .B(n3563), .Z(n3473) );
  IV U1446 ( .A(n3583), .Z(n3563) );
  AN2 U1447 ( .A(n3584), .B(n3585), .Z(n3583) );
  AN2 U1448 ( .A(n262), .B(n195), .Z(n3585) );
  AN2 U1449 ( .A(n461), .B(n328), .Z(n3584) );
  IV U1450 ( .A(n3586), .Z(n3558) );
  AN2 U1451 ( .A(n3587), .B(n3588), .Z(n3586) );
  AN2 U1452 ( .A(n229), .B(n159), .Z(n3588) );
  AN2 U1453 ( .A(n428), .B(n295), .Z(n3587) );
  OR2 U1454 ( .A(n3499), .B(n3576), .Z(n3582) );
  OR2 U1455 ( .A(n3498), .B(n3493), .Z(n3576) );
  IV U1456 ( .A(n616), .Z(n3493) );
  IV U1457 ( .A(n176), .Z(n3498) );
  IV U1458 ( .A(n191), .Z(n3499) );
  AN2 U1459 ( .A(n3589), .B(n3506), .Z(n3579) );
  IV U1460 ( .A(n615), .Z(n3506) );
  OR2 U1461 ( .A(n3469), .B(n3501), .Z(n3589) );
  IV U1462 ( .A(n619), .Z(n3501) );
  OR2 U1463 ( .A(n3486), .B(n3540), .Z(n3469) );
  IV U1464 ( .A(n3590), .Z(n3540) );
  AN2 U1465 ( .A(n3591), .B(n3592), .Z(n3590) );
  AN2 U1466 ( .A(n572), .B(n580), .Z(n3592) );
  AN2 U1467 ( .A(n593), .B(n577), .Z(n3591) );
  IV U1468 ( .A(n3593), .Z(n3486) );
  AN2 U1469 ( .A(n627), .B(n622), .Z(n3593) );
  AN2 U1470 ( .A(n678), .B(n3594), .Z(n3520) );
  IV U1471 ( .A(n48), .Z(n3518) );
  OR2 U1472 ( .A(n3595), .B(n2447), .Z(U50_Z_7) );
  AN2 U1473 ( .A(U50_DATA1_7), .B(U50_CONTROL1), .Z(n3595) );
  OR2 U1474 ( .A(n3596), .B(n3597), .Z(U50_Z_6) );
  OR2 U1475 ( .A(n2451), .B(n2448), .Z(n3597) );
  AN2 U1476 ( .A(U50_DATA1_6), .B(U50_CONTROL1), .Z(n3596) );
  OR2 U1477 ( .A(n3598), .B(n3599), .Z(U50_Z_5) );
  OR2 U1478 ( .A(n2455), .B(n2452), .Z(n3599) );
  AN2 U1479 ( .A(U50_DATA1_5), .B(U50_CONTROL1), .Z(n3598) );
  OR2 U1480 ( .A(n3600), .B(n2457), .Z(U50_Z_4) );
  AN2 U1481 ( .A(U50_DATA1_4), .B(U50_CONTROL1), .Z(n3600) );
  OR2 U1482 ( .A(n3601), .B(n3602), .Z(U50_Z_3) );
  OR2 U1483 ( .A(n2461), .B(n2458), .Z(n3602) );
  AN2 U1484 ( .A(U50_CONTROL1), .B(U50_DATA1_3), .Z(n3601) );
  OR2 U1485 ( .A(n3603), .B(n3604), .Z(U50_Z_2) );
  OR2 U1486 ( .A(n2465), .B(n2462), .Z(n3604) );
  AN2 U1487 ( .A(U50_CONTROL1), .B(U50_DATA1_2), .Z(n3603) );
  OR2 U1488 ( .A(n3605), .B(n3606), .Z(U50_Z_1) );
  OR2 U1489 ( .A(n2469), .B(n2466), .Z(n3606) );
  AN2 U1490 ( .A(U50_CONTROL1), .B(U50_DATA1_1), .Z(n3605) );
  OR2 U1491 ( .A(n3607), .B(n3608), .Z(U50_Z_0) );
  OR2 U1492 ( .A(n2473), .B(n2470), .Z(n3608) );
  AN2 U1493 ( .A(U50_CONTROL1), .B(U50_DATA1_0), .Z(n3607) );
  OR2 U1494 ( .A(n3609), .B(n3610), .Z(U5_Z_9) );
  AN2 U1495 ( .A(U5_DATA1_9), .B(n3611), .Z(n3609) );
  AN2 U1496 ( .A(U5_DATA1_8), .B(n3611), .Z(U5_Z_8) );
  OR2 U1497 ( .A(n3612), .B(n3613), .Z(U5_Z_7) );
  AN2 U1498 ( .A(U5_DATA1_7), .B(n3611), .Z(n3612) );
  OR2 U1499 ( .A(n3614), .B(n28), .Z(U5_Z_6) );
  AN2 U1500 ( .A(U5_DATA1_6), .B(n3611), .Z(n3614) );
  OR2 U1501 ( .A(n3615), .B(n3613), .Z(U5_Z_5) );
  AN2 U1502 ( .A(U5_DATA1_5), .B(n3611), .Z(n3615) );
  OR2 U1503 ( .A(n3616), .B(n28), .Z(U5_Z_4) );
  AN2 U1504 ( .A(U5_DATA1_4), .B(n3611), .Z(n3616) );
  OR2 U1505 ( .A(n3617), .B(n3613), .Z(U5_Z_3) );
  OR2 U1506 ( .A(n3610), .B(n28), .Z(n3613) );
  AN2 U1507 ( .A(U5_DATA1_3), .B(n3611), .Z(n3617) );
  AN2 U1508 ( .A(U5_DATA1_2), .B(n3611), .Z(U5_Z_2) );
  OR2 U1509 ( .A(n3618), .B(n3610), .Z(U5_Z_1) );
  AN2 U1510 ( .A(n3619), .B(n[2079]), .Z(n3610) );
  AN2 U1511 ( .A(U5_DATA1_1), .B(n3611), .Z(n3618) );
  AN2 U1512 ( .A(U5_DATA1_0), .B(n3611), .Z(U5_Z_0) );
  AN2 U1513 ( .A(n3619), .B(n3517), .Z(n3611) );
  IV U1514 ( .A(n[2079]), .Z(n3517) );
  IV U1515 ( .A(n[2080]), .Z(n3619) );
  OR2 U1516 ( .A(n3620), .B(n2484), .Z(U4_Z_3) );
  AN2 U1517 ( .A(U4_DATA2_3), .B(link_up_loc), .Z(n3620) );
  OR2 U1518 ( .A(n3621), .B(n2486), .Z(U4_Z_2) );
  AN2 U1519 ( .A(U4_DATA2_2), .B(link_up_loc), .Z(n3621) );
  OR2 U1520 ( .A(n3622), .B(n2488), .Z(U4_Z_1) );
  AN2 U1521 ( .A(U4_DATA2_1), .B(link_up_loc), .Z(n3622) );
  OR2 U1522 ( .A(n3623), .B(n2490), .Z(U4_Z_0) );
  AN2 U1523 ( .A(link_up_loc), .B(U4_DATA2_0), .Z(n3623) );
  OR2 U1524 ( .A(n3624), .B(n3625), .Z(U20_Z_9) );
  AN2 U1525 ( .A(n3626), .B(n3528), .Z(n3625) );
  OR2 U1526 ( .A(n3627), .B(n3628), .Z(n3626) );
  OR2 U1527 ( .A(n3629), .B(n3630), .Z(n3628) );
  OR2 U1528 ( .A(n3631), .B(n3632), .Z(n3630) );
  OR2 U1529 ( .A(n3633), .B(n3634), .Z(n3632) );
  AN2 U1530 ( .A(U47_DATA121_0), .B(n3635), .Z(n3634) );
  AN2 U1531 ( .A(n3636), .B(n3531), .Z(n3633) );
  OR2 U1532 ( .A(n3637), .B(n3638), .Z(n3629) );
  OR2 U1533 ( .A(n3639), .B(n3640), .Z(n3638) );
  OR2 U1534 ( .A(n3641), .B(n3642), .Z(n3627) );
  OR2 U1535 ( .A(n3643), .B(n3644), .Z(n3642) );
  AN2 U1536 ( .A(n3645), .B(n3646), .Z(n3643) );
  OR2 U1537 ( .A(n3647), .B(n3648), .Z(n3641) );
  OR2 U1538 ( .A(n1893), .B(n3649), .Z(n3648) );
  AN2 U1539 ( .A(n3650), .B(n3651), .Z(n3647) );
  AN2 U1540 ( .A(n2112), .B(n3652), .Z(n3624) );
  OR2 U1541 ( .A(n1919), .B(n3653), .Z(n3652) );
  OR2 U1542 ( .A(n3654), .B(n3655), .Z(n3653) );
  AN2 U1543 ( .A(U47_DATA121_0), .B(n3656), .Z(n3655) );
  OR2 U1544 ( .A(n3657), .B(n3658), .Z(n3656) );
  AN2 U1545 ( .A(n3659), .B(n3531), .Z(n3654) );
  OR2 U1546 ( .A(n3660), .B(n3661), .Z(n3659) );
  OR2 U1547 ( .A(n3662), .B(n2311), .Z(n3661) );
  OR2 U1548 ( .A(n3663), .B(n3664), .Z(U20_Z_8) );
  OR2 U1549 ( .A(n3665), .B(n3666), .Z(n3664) );
  AN2 U1550 ( .A(n3667), .B(n3528), .Z(n3666) );
  OR2 U1551 ( .A(n3668), .B(n3669), .Z(n3667) );
  OR2 U1552 ( .A(n3670), .B(n3671), .Z(n3669) );
  OR2 U1553 ( .A(n3672), .B(n3673), .Z(n3671) );
  OR2 U1554 ( .A(n3674), .B(n3675), .Z(n3673) );
  AN2 U1555 ( .A(U47_DATA121_0), .B(n3676), .Z(n3675) );
  AN2 U1556 ( .A(n3677), .B(n3531), .Z(n3674) );
  OR2 U1557 ( .A(n3678), .B(n3679), .Z(n3670) );
  OR2 U1558 ( .A(n3680), .B(n3681), .Z(n3679) );
  OR2 U1559 ( .A(n3682), .B(n3683), .Z(n3668) );
  OR2 U1560 ( .A(n3684), .B(n3685), .Z(n3683) );
  OR2 U1561 ( .A(n3686), .B(n3687), .Z(n3685) );
  AN2 U1562 ( .A(n3688), .B(n3651), .Z(n3687) );
  AN2 U1563 ( .A(n3689), .B(n3645), .Z(n3684) );
  OR2 U1564 ( .A(n3690), .B(n3691), .Z(n3682) );
  OR2 U1565 ( .A(n1855), .B(n3448), .Z(n3691) );
  AN2 U1566 ( .A(n3524), .B(n3692), .Z(n3665) );
  OR2 U1567 ( .A(n3693), .B(n3694), .Z(n3692) );
  AN2 U1568 ( .A(n3594), .B(n3695), .Z(n3663) );
  OR2 U1569 ( .A(n3696), .B(n3697), .Z(U20_Z_7) );
  OR2 U1570 ( .A(n3698), .B(n3699), .Z(n3697) );
  AN2 U1571 ( .A(n3524), .B(n3700), .Z(n3699) );
  OR2 U1572 ( .A(n3695), .B(n3701), .Z(n3700) );
  OR2 U1573 ( .A(n3657), .B(n3694), .Z(n3701) );
  AN2 U1574 ( .A(n3662), .B(n3594), .Z(n3698) );
  OR2 U1575 ( .A(n3702), .B(n3703), .Z(n3696) );
  AN2 U1576 ( .A(n3704), .B(n3528), .Z(n3703) );
  OR2 U1577 ( .A(n3705), .B(n3706), .Z(n3704) );
  OR2 U1578 ( .A(n3707), .B(n3708), .Z(n3706) );
  OR2 U1579 ( .A(n3709), .B(n3710), .Z(n3708) );
  OR2 U1580 ( .A(n3711), .B(n3712), .Z(n3710) );
  AN2 U1581 ( .A(U47_DATA121_0), .B(n3713), .Z(n3712) );
  AN2 U1582 ( .A(n3714), .B(n3531), .Z(n3711) );
  OR2 U1583 ( .A(n3715), .B(n3716), .Z(n3707) );
  OR2 U1584 ( .A(n3640), .B(n3717), .Z(n3716) );
  OR2 U1585 ( .A(n3718), .B(n3719), .Z(n3705) );
  OR2 U1586 ( .A(n3720), .B(n3639), .Z(n3719) );
  OR2 U1587 ( .A(n3721), .B(n3722), .Z(n3639) );
  OR2 U1588 ( .A(n3723), .B(n3724), .Z(n3722) );
  AN2 U1589 ( .A(n3725), .B(n3651), .Z(n3724) );
  AN2 U1590 ( .A(n3726), .B(n3531), .Z(n3723) );
  AN2 U1591 ( .A(n3645), .B(n3727), .Z(n3721) );
  OR2 U1592 ( .A(n3728), .B(n3729), .Z(n3718) );
  OR2 U1593 ( .A(n1836), .B(n3730), .Z(n3729) );
  AN2 U1594 ( .A(n3731), .B(n3651), .Z(n3730) );
  AN2 U1595 ( .A(n3645), .B(n3732), .Z(n3728) );
  OR2 U1596 ( .A(n3733), .B(n3734), .Z(U20_Z_6) );
  OR2 U1597 ( .A(n3735), .B(n3736), .Z(n3734) );
  AN2 U1598 ( .A(n3594), .B(n3694), .Z(n3736) );
  OR2 U1599 ( .A(n3737), .B(n2312), .Z(n3694) );
  AN2 U1600 ( .A(n3738), .B(n3739), .Z(n3737) );
  AN2 U1601 ( .A(n3524), .B(n3740), .Z(n3735) );
  OR2 U1602 ( .A(n3693), .B(n3695), .Z(n3740) );
  OR2 U1603 ( .A(n3741), .B(n3742), .Z(n3695) );
  OR2 U1604 ( .A(n3743), .B(n2311), .Z(n3742) );
  AN2 U1605 ( .A(n3738), .B(n3744), .Z(n3741) );
  AN2 U1606 ( .A(n3745), .B(n3528), .Z(n3733) );
  OR2 U1607 ( .A(n3746), .B(n3747), .Z(n3745) );
  OR2 U1608 ( .A(n3748), .B(n3749), .Z(n3747) );
  OR2 U1609 ( .A(n3750), .B(n3751), .Z(n3749) );
  OR2 U1610 ( .A(n3752), .B(n3753), .Z(n3751) );
  AN2 U1611 ( .A(n3676), .B(n3531), .Z(n3753) );
  OR2 U1612 ( .A(n3754), .B(n3755), .Z(n3676) );
  OR2 U1613 ( .A(n3756), .B(n3714), .Z(n3755) );
  AN2 U1614 ( .A(U47_DATA121_0), .B(n3677), .Z(n3752) );
  OR2 U1615 ( .A(n3726), .B(n3757), .Z(n3677) );
  OR2 U1616 ( .A(n3758), .B(n3759), .Z(n3757) );
  OR2 U1617 ( .A(n3760), .B(n3761), .Z(n3726) );
  OR2 U1618 ( .A(n3762), .B(n3763), .Z(n3748) );
  OR2 U1619 ( .A(n3640), .B(n3678), .Z(n3763) );
  OR2 U1620 ( .A(n3764), .B(n3765), .Z(n3678) );
  OR2 U1621 ( .A(n3766), .B(n3767), .Z(n3765) );
  OR2 U1622 ( .A(n3768), .B(n3769), .Z(n3767) );
  AN2 U1623 ( .A(n3770), .B(n3531), .Z(n3769) );
  OR2 U1624 ( .A(n3771), .B(n3772), .Z(n3770) );
  OR2 U1625 ( .A(n3773), .B(n3774), .Z(n3772) );
  OR2 U1626 ( .A(n3775), .B(n3776), .Z(n3771) );
  OR2 U1627 ( .A(n3777), .B(n3778), .Z(n3776) );
  AN2 U1628 ( .A(U47_DATA121_0), .B(n3779), .Z(n3768) );
  OR2 U1629 ( .A(n3780), .B(n3781), .Z(n3764) );
  OR2 U1630 ( .A(n3637), .B(n3717), .Z(n3781) );
  OR2 U1631 ( .A(n3782), .B(n3783), .Z(n3717) );
  OR2 U1632 ( .A(n3445), .B(n3784), .Z(n3783) );
  AN2 U1633 ( .A(n3785), .B(n3731), .Z(n3784) );
  AN2 U1634 ( .A(n3786), .B(n3787), .Z(n3782) );
  OR2 U1635 ( .A(n3788), .B(n3789), .Z(n3637) );
  AN2 U1636 ( .A(n3785), .B(n3650), .Z(n3789) );
  AN2 U1637 ( .A(n3790), .B(n3791), .Z(n3788) );
  OR2 U1638 ( .A(n3792), .B(n3793), .Z(n3640) );
  OR2 U1639 ( .A(n3449), .B(n3794), .Z(n3793) );
  AN2 U1640 ( .A(n3785), .B(n3725), .Z(n3794) );
  AN2 U1641 ( .A(n3786), .B(n3795), .Z(n3792) );
  OR2 U1642 ( .A(n3796), .B(n3797), .Z(n3746) );
  OR2 U1643 ( .A(n3798), .B(n3799), .Z(n3797) );
  OR2 U1644 ( .A(n3800), .B(n3801), .Z(n3796) );
  OR2 U1645 ( .A(n3802), .B(n3803), .Z(U20_Z_5) );
  OR2 U1646 ( .A(n3804), .B(n3805), .Z(n3803) );
  AN2 U1647 ( .A(n2312), .B(n3524), .Z(n3804) );
  OR2 U1648 ( .A(n3806), .B(n3807), .Z(n3802) );
  AN2 U1649 ( .A(n2311), .B(n3594), .Z(n3807) );
  AN2 U1650 ( .A(n3808), .B(n3528), .Z(n3806) );
  OR2 U1651 ( .A(n3809), .B(n3810), .Z(n3808) );
  OR2 U1652 ( .A(n3811), .B(n3812), .Z(n3810) );
  OR2 U1653 ( .A(n3709), .B(n3813), .Z(n3812) );
  OR2 U1654 ( .A(n3814), .B(n3815), .Z(n3813) );
  AN2 U1655 ( .A(n3816), .B(n3531), .Z(n3815) );
  OR2 U1656 ( .A(n3817), .B(n3713), .Z(n3816) );
  OR2 U1657 ( .A(n3818), .B(n3819), .Z(n3713) );
  OR2 U1658 ( .A(n3778), .B(n3775), .Z(n3819) );
  OR2 U1659 ( .A(n3756), .B(n3759), .Z(n3818) );
  AN2 U1660 ( .A(U47_DATA121_0), .B(n3820), .Z(n3814) );
  OR2 U1661 ( .A(n3761), .B(n3821), .Z(n3820) );
  OR2 U1662 ( .A(n3714), .B(n3822), .Z(n3821) );
  OR2 U1663 ( .A(n3823), .B(n3824), .Z(n3709) );
  OR2 U1664 ( .A(n3825), .B(n3826), .Z(n3824) );
  OR2 U1665 ( .A(n3686), .B(n3762), .Z(n3826) );
  OR2 U1666 ( .A(n3827), .B(n3828), .Z(n3762) );
  AN2 U1667 ( .A(n3645), .B(n3829), .Z(n3828) );
  AN2 U1668 ( .A(n3830), .B(n3831), .Z(n3827) );
  AN2 U1669 ( .A(n3832), .B(n3830), .Z(n3686) );
  OR2 U1670 ( .A(n3833), .B(n3834), .Z(n3825) );
  AN2 U1671 ( .A(n3835), .B(n3531), .Z(n3834) );
  OR2 U1672 ( .A(n3836), .B(n3837), .Z(n3835) );
  OR2 U1673 ( .A(n3754), .B(n3774), .Z(n3837) );
  OR2 U1674 ( .A(n3758), .B(n3779), .Z(n3836) );
  AN2 U1675 ( .A(U47_DATA121_0), .B(n3777), .Z(n3833) );
  OR2 U1676 ( .A(n3838), .B(n3839), .Z(n3823) );
  OR2 U1677 ( .A(n3840), .B(n3649), .Z(n3839) );
  AN2 U1678 ( .A(n3841), .B(n3830), .Z(n3649) );
  OR2 U1679 ( .A(n3451), .B(n3444), .Z(n3838) );
  OR2 U1680 ( .A(n3780), .B(n3842), .Z(n3811) );
  OR2 U1681 ( .A(n3843), .B(n3644), .Z(n3842) );
  OR2 U1682 ( .A(n3799), .B(n3844), .Z(n3644) );
  OR2 U1683 ( .A(n3845), .B(n3681), .Z(n3844) );
  OR2 U1684 ( .A(n3846), .B(n3847), .Z(n3681) );
  AN2 U1685 ( .A(n3830), .B(n3848), .Z(n3846) );
  AN2 U1686 ( .A(U47_DATA121_0), .B(n3773), .Z(n3845) );
  OR2 U1687 ( .A(n3849), .B(n3850), .Z(n3799) );
  AN2 U1688 ( .A(n3645), .B(n3851), .Z(n3850) );
  AN2 U1689 ( .A(n3830), .B(n3852), .Z(n3849) );
  OR2 U1690 ( .A(n3853), .B(n3854), .Z(n3780) );
  AN2 U1691 ( .A(n3645), .B(n3855), .Z(n3854) );
  AN2 U1692 ( .A(n3830), .B(n3856), .Z(n3853) );
  OR2 U1693 ( .A(n3857), .B(n3858), .Z(n3809) );
  OR2 U1694 ( .A(n3690), .B(n3859), .Z(n3858) );
  OR2 U1695 ( .A(n3447), .B(n3860), .Z(n3859) );
  OR2 U1696 ( .A(n3448), .B(n3801), .Z(n3857) );
  OR2 U1697 ( .A(n1730), .B(n3450), .Z(n3801) );
  OR2 U1698 ( .A(n3861), .B(n3862), .Z(U20_Z_4) );
  OR2 U1699 ( .A(n3863), .B(n3864), .Z(n3862) );
  AN2 U1700 ( .A(n3524), .B(n3865), .Z(n3863) );
  OR2 U1701 ( .A(n2311), .B(n3658), .Z(n3865) );
  OR2 U1702 ( .A(n3743), .B(n2312), .Z(n3658) );
  OR2 U1703 ( .A(n3866), .B(n3867), .Z(n3861) );
  AN2 U1704 ( .A(n3868), .B(n3528), .Z(n3867) );
  OR2 U1705 ( .A(n3869), .B(n3870), .Z(n3868) );
  OR2 U1706 ( .A(n3871), .B(n3872), .Z(n3870) );
  OR2 U1707 ( .A(n3715), .B(n3873), .Z(n3872) );
  OR2 U1708 ( .A(n3874), .B(n3875), .Z(n3873) );
  AN2 U1709 ( .A(n3876), .B(n3531), .Z(n3875) );
  OR2 U1710 ( .A(n3761), .B(n3635), .Z(n3876) );
  OR2 U1711 ( .A(n3758), .B(n3778), .Z(n3635) );
  OR2 U1712 ( .A(n3877), .B(n3878), .Z(n3778) );
  AN2 U1713 ( .A(n3879), .B(n3880), .Z(n3878) );
  AN2 U1714 ( .A(n3790), .B(n3881), .Z(n3877) );
  AN2 U1715 ( .A(n3882), .B(n3883), .Z(n3758) );
  OR2 U1716 ( .A(n3830), .B(n3884), .Z(n3883) );
  OR2 U1717 ( .A(n3885), .B(n3886), .Z(n3761) );
  AN2 U1718 ( .A(n3887), .B(n3888), .Z(n3886) );
  AN2 U1719 ( .A(n3889), .B(n3890), .Z(n3885) );
  AN2 U1720 ( .A(U47_DATA121_0), .B(n3891), .Z(n3874) );
  OR2 U1721 ( .A(n3760), .B(n3636), .Z(n3891) );
  OR2 U1722 ( .A(n3775), .B(n3754), .Z(n3636) );
  OR2 U1723 ( .A(n3892), .B(n3893), .Z(n3754) );
  AN2 U1724 ( .A(n3830), .B(n3725), .Z(n3893) );
  AN2 U1725 ( .A(n3894), .B(n3795), .Z(n3892) );
  OR2 U1726 ( .A(n3895), .B(n3896), .Z(n3775) );
  AN2 U1727 ( .A(n3830), .B(n3650), .Z(n3896) );
  AN2 U1728 ( .A(n3894), .B(n3791), .Z(n3895) );
  OR2 U1729 ( .A(n3817), .B(n3822), .Z(n3760) );
  OR2 U1730 ( .A(n3897), .B(n3898), .Z(n3822) );
  AN2 U1731 ( .A(n3879), .B(n3899), .Z(n3898) );
  AN2 U1732 ( .A(n3790), .B(n3900), .Z(n3897) );
  OR2 U1733 ( .A(n3901), .B(n3902), .Z(n3817) );
  AN2 U1734 ( .A(n3830), .B(n3899), .Z(n3902) );
  AN2 U1735 ( .A(n3894), .B(n3900), .Z(n3901) );
  OR2 U1736 ( .A(n3903), .B(n3904), .Z(n3715) );
  OR2 U1737 ( .A(n3672), .B(n3750), .Z(n3904) );
  OR2 U1738 ( .A(n3905), .B(n3906), .Z(n3750) );
  AN2 U1739 ( .A(n3785), .B(n3831), .Z(n3906) );
  AN2 U1740 ( .A(n3790), .B(n3829), .Z(n3905) );
  OR2 U1741 ( .A(n3907), .B(n3908), .Z(n3672) );
  AN2 U1742 ( .A(n3879), .B(n3832), .Z(n3908) );
  AN2 U1743 ( .A(n3790), .B(n3732), .Z(n3907) );
  OR2 U1744 ( .A(n3909), .B(n3910), .Z(n3903) );
  OR2 U1745 ( .A(n3911), .B(n3912), .Z(n3910) );
  AN2 U1746 ( .A(n3831), .B(n3651), .Z(n3912) );
  AN2 U1747 ( .A(n3773), .B(n3531), .Z(n3911) );
  OR2 U1748 ( .A(n3913), .B(n3914), .Z(n3773) );
  AN2 U1749 ( .A(n3915), .B(n3916), .Z(n3914) );
  AN2 U1750 ( .A(n3889), .B(n3917), .Z(n3913) );
  AN2 U1751 ( .A(n3645), .B(n3918), .Z(n3909) );
  OR2 U1752 ( .A(n3631), .B(n3766), .Z(n3871) );
  OR2 U1753 ( .A(n3919), .B(n3920), .Z(n3766) );
  AN2 U1754 ( .A(n3785), .B(n3856), .Z(n3920) );
  AN2 U1755 ( .A(n3790), .B(n3855), .Z(n3919) );
  OR2 U1756 ( .A(n3786), .B(n3887), .Z(n3790) );
  OR2 U1757 ( .A(n3921), .B(n3922), .Z(n3631) );
  OR2 U1758 ( .A(n3843), .B(n3923), .Z(n3922) );
  OR2 U1759 ( .A(n3924), .B(n3925), .Z(n3923) );
  AN2 U1760 ( .A(n3926), .B(n3531), .Z(n3925) );
  OR2 U1761 ( .A(n3927), .B(n3928), .Z(n3926) );
  OR2 U1762 ( .A(n3759), .B(n3779), .Z(n3928) );
  OR2 U1763 ( .A(n3929), .B(n3930), .Z(n3779) );
  OR2 U1764 ( .A(n3931), .B(n3932), .Z(n3930) );
  AN2 U1765 ( .A(n3645), .B(n3881), .Z(n3932) );
  AN2 U1766 ( .A(n3830), .B(n3880), .Z(n3931) );
  OR2 U1767 ( .A(n3933), .B(n3934), .Z(n3759) );
  AN2 U1768 ( .A(n3830), .B(n3890), .Z(n3934) );
  AN2 U1769 ( .A(n3894), .B(n3888), .Z(n3933) );
  OR2 U1770 ( .A(n3714), .B(n3935), .Z(n3927) );
  OR2 U1771 ( .A(n3777), .B(n3756), .Z(n3935) );
  OR2 U1772 ( .A(n3936), .B(n3937), .Z(n3756) );
  AN2 U1773 ( .A(n3938), .B(n3882), .Z(n3936) );
  OR2 U1774 ( .A(n3939), .B(n3940), .Z(n3938) );
  OR2 U1775 ( .A(n3786), .B(n3915), .Z(n3940) );
  OR2 U1776 ( .A(n3941), .B(n3651), .Z(n3939) );
  OR2 U1777 ( .A(n3942), .B(n3943), .Z(n3777) );
  AN2 U1778 ( .A(n3887), .B(n3918), .Z(n3943) );
  AN2 U1779 ( .A(n3889), .B(n3944), .Z(n3942) );
  OR2 U1780 ( .A(n3945), .B(n3946), .Z(n3714) );
  AN2 U1781 ( .A(n3887), .B(n3947), .Z(n3946) );
  AN2 U1782 ( .A(n3889), .B(n3948), .Z(n3945) );
  AN2 U1783 ( .A(U47_DATA121_0), .B(n3774), .Z(n3924) );
  OR2 U1784 ( .A(n3949), .B(n3950), .Z(n3774) );
  AN2 U1785 ( .A(n3830), .B(n3731), .Z(n3950) );
  AN2 U1786 ( .A(n3894), .B(n3787), .Z(n3949) );
  OR2 U1787 ( .A(n3951), .B(n3645), .Z(n3894) );
  OR2 U1788 ( .A(n3952), .B(n3953), .Z(n3843) );
  AN2 U1789 ( .A(n3830), .B(n3917), .Z(n3953) );
  AN2 U1790 ( .A(n3884), .B(n3916), .Z(n3952) );
  OR2 U1791 ( .A(n3954), .B(n3951), .Z(n3884) );
  OR2 U1792 ( .A(n3680), .B(n3955), .Z(n3921) );
  OR2 U1793 ( .A(n3720), .B(n3798), .Z(n3955) );
  OR2 U1794 ( .A(n3956), .B(n3957), .Z(n3798) );
  OR2 U1795 ( .A(n3958), .B(n3959), .Z(n3957) );
  AN2 U1796 ( .A(n3786), .B(n3960), .Z(n3959) );
  AN2 U1797 ( .A(n3879), .B(n3852), .Z(n3958) );
  AN2 U1798 ( .A(n3887), .B(n3851), .Z(n3956) );
  OR2 U1799 ( .A(n3961), .B(n3962), .Z(n3720) );
  OR2 U1800 ( .A(n3963), .B(n3964), .Z(n3962) );
  AN2 U1801 ( .A(n3786), .B(n3965), .Z(n3964) );
  AN2 U1802 ( .A(n3879), .B(n3841), .Z(n3963) );
  AN2 U1803 ( .A(n3887), .B(n3727), .Z(n3961) );
  OR2 U1804 ( .A(n3966), .B(n3967), .Z(n3680) );
  AN2 U1805 ( .A(n3887), .B(n3646), .Z(n3967) );
  AN2 U1806 ( .A(n3889), .B(n3848), .Z(n3966) );
  OR2 U1807 ( .A(n3879), .B(n3786), .Z(n3889) );
  OR2 U1808 ( .A(n3785), .B(n3651), .Z(n3879) );
  OR2 U1809 ( .A(n3941), .B(n3968), .Z(n3785) );
  OR2 U1810 ( .A(n3969), .B(n3970), .Z(n3941) );
  OR2 U1811 ( .A(n3971), .B(n3972), .Z(n3970) );
  OR2 U1812 ( .A(n3973), .B(n3974), .Z(n3969) );
  OR2 U1813 ( .A(n3975), .B(n3976), .Z(n3869) );
  OR2 U1814 ( .A(n3977), .B(n3978), .Z(n3976) );
  AN2 U1815 ( .A(n3645), .B(n3947), .Z(n3978) );
  AN2 U1816 ( .A(n3856), .B(n3651), .Z(n3977) );
  OR2 U1817 ( .A(n3840), .B(n3979), .Z(n3975) );
  OR2 U1818 ( .A(n1643), .B(n3690), .Z(n3979) );
  AN2 U1819 ( .A(n3948), .B(n3830), .Z(n3690) );
  AN2 U1820 ( .A(n3944), .B(n3830), .Z(n3840) );
  OR2 U1821 ( .A(n3980), .B(n3981), .Z(n3830) );
  OR2 U1822 ( .A(n3982), .B(n3983), .Z(n3981) );
  OR2 U1823 ( .A(n3984), .B(n3985), .Z(n3983) );
  OR2 U1824 ( .A(n3986), .B(n3987), .Z(n3980) );
  OR2 U1825 ( .A(n3988), .B(n3989), .Z(n3987) );
  AN2 U1826 ( .A(n2318), .B(n2112), .Z(n3866) );
  OR2 U1827 ( .A(n3990), .B(n3805), .Z(U20_Z_3) );
  OR2 U1828 ( .A(n3991), .B(n3992), .Z(n3805) );
  AN2 U1829 ( .A(n2316), .B(n2112), .Z(n3992) );
  AN2 U1830 ( .A(n3993), .B(n3744), .Z(n2316) );
  AN2 U1831 ( .A(n3524), .B(n3994), .Z(n3991) );
  AN2 U1832 ( .A(n3995), .B(n3528), .Z(n3990) );
  OR2 U1833 ( .A(n3996), .B(n3997), .Z(n3995) );
  OR2 U1834 ( .A(n3998), .B(n3999), .Z(n3997) );
  OR2 U1835 ( .A(n4000), .B(n4001), .Z(n3999) );
  OR2 U1836 ( .A(n4002), .B(n4003), .Z(n3998) );
  AN2 U1837 ( .A(n4004), .B(n3531), .Z(n4002) );
  OR2 U1838 ( .A(n4005), .B(n4006), .Z(n3996) );
  OR2 U1839 ( .A(n1661), .B(n4007), .Z(n4006) );
  OR2 U1840 ( .A(n4008), .B(n4009), .Z(U20_Z_2) );
  OR2 U1841 ( .A(n4010), .B(n4011), .Z(n4009) );
  AN2 U1842 ( .A(n2112), .B(n4012), .Z(n4011) );
  OR2 U1843 ( .A(n2311), .B(n4013), .Z(n4012) );
  OR2 U1844 ( .A(n2318), .B(n2312), .Z(n4013) );
  AN2 U1845 ( .A(n4014), .B(n3739), .Z(n2312) );
  AN2 U1846 ( .A(n3738), .B(n4015), .Z(n2318) );
  AN2 U1847 ( .A(n3993), .B(n3739), .Z(n2311) );
  IV U1848 ( .A(n1615), .Z(n3993) );
  AN2 U1849 ( .A(n4016), .B(n3528), .Z(n4010) );
  OR2 U1850 ( .A(n4017), .B(n4018), .Z(n4016) );
  OR2 U1851 ( .A(n4019), .B(n4020), .Z(n4018) );
  OR2 U1852 ( .A(n4021), .B(n4022), .Z(n4020) );
  AN2 U1853 ( .A(U47_DATA121_0), .B(n4023), .Z(n4022) );
  OR2 U1854 ( .A(n4024), .B(n4004), .Z(n4023) );
  AN2 U1855 ( .A(n4025), .B(n3531), .Z(n4021) );
  OR2 U1856 ( .A(n4026), .B(n4005), .Z(n4017) );
  OR2 U1857 ( .A(n4027), .B(n4028), .Z(n4005) );
  AN2 U1858 ( .A(n4029), .B(n3531), .Z(n4028) );
  OR2 U1859 ( .A(n4030), .B(n4031), .Z(n4029) );
  AN2 U1860 ( .A(U47_DATA121_0), .B(n4032), .Z(n4027) );
  OR2 U1861 ( .A(n4033), .B(n4034), .Z(U20_Z_1) );
  OR2 U1862 ( .A(n4035), .B(n3864), .Z(n4034) );
  AN2 U1863 ( .A(n3594), .B(n4036), .Z(n3864) );
  AN2 U1864 ( .A(n3743), .B(n3524), .Z(n4035) );
  AN2 U1865 ( .A(n3531), .B(n2112), .Z(n3524) );
  OR2 U1866 ( .A(n3702), .B(n4037), .Z(n4033) );
  AN2 U1867 ( .A(n4038), .B(n3528), .Z(n4037) );
  OR2 U1868 ( .A(n4039), .B(n4040), .Z(n4038) );
  OR2 U1869 ( .A(n4041), .B(n4042), .Z(n4040) );
  OR2 U1870 ( .A(n4043), .B(n4044), .Z(n4042) );
  AN2 U1871 ( .A(U47_DATA121_0), .B(n4031), .Z(n4044) );
  AN2 U1872 ( .A(n4045), .B(n3531), .Z(n4043) );
  OR2 U1873 ( .A(n4000), .B(n4026), .Z(n4039) );
  OR2 U1874 ( .A(n4046), .B(n4047), .Z(n4026) );
  OR2 U1875 ( .A(n4048), .B(n4049), .Z(n4047) );
  AN2 U1876 ( .A(n4050), .B(n3786), .Z(n4049) );
  IV U1877 ( .A(n1414), .Z(n3786) );
  OR2 U1878 ( .A(n4051), .B(n4052), .Z(n4050) );
  OR2 U1879 ( .A(n4053), .B(n4054), .Z(n4052) );
  OR2 U1880 ( .A(n3960), .B(n4055), .Z(n4054) );
  OR2 U1881 ( .A(n3829), .B(n3965), .Z(n4055) );
  IV U1882 ( .A(n1425), .Z(n3965) );
  IV U1883 ( .A(n1434), .Z(n3960) );
  OR2 U1884 ( .A(n3855), .B(n4056), .Z(n4053) );
  OR2 U1885 ( .A(n3900), .B(n3881), .Z(n4056) );
  OR2 U1886 ( .A(n4057), .B(n4058), .Z(n4051) );
  OR2 U1887 ( .A(n4059), .B(n4060), .Z(n4058) );
  OR2 U1888 ( .A(n3882), .B(n4061), .Z(n4060) );
  OR2 U1889 ( .A(n3890), .B(n4062), .Z(n4057) );
  OR2 U1890 ( .A(n3732), .B(n3848), .Z(n4062) );
  AN2 U1891 ( .A(n4063), .B(n3531), .Z(n4048) );
  OR2 U1892 ( .A(n4064), .B(n4065), .Z(n4063) );
  OR2 U1893 ( .A(n4007), .B(n4066), .Z(n4065) );
  OR2 U1894 ( .A(n3444), .B(n4067), .Z(n4066) );
  AN2 U1895 ( .A(n3951), .B(n3918), .Z(n3444) );
  AN2 U1896 ( .A(n3887), .B(n3791), .Z(n4007) );
  OR2 U1897 ( .A(n3445), .B(n4068), .Z(n4064) );
  OR2 U1898 ( .A(n3449), .B(n3448), .Z(n4068) );
  AN2 U1899 ( .A(n3951), .B(n3947), .Z(n3448) );
  AN2 U1900 ( .A(n3795), .B(n3887), .Z(n3449) );
  AN2 U1901 ( .A(n3787), .B(n3887), .Z(n3445) );
  OR2 U1902 ( .A(n4069), .B(n4070), .Z(n4046) );
  OR2 U1903 ( .A(n3860), .B(n4071), .Z(n4070) );
  AN2 U1904 ( .A(n4072), .B(n3645), .Z(n4071) );
  OR2 U1905 ( .A(n4073), .B(n4074), .Z(n4072) );
  OR2 U1906 ( .A(n4075), .B(n3881), .Z(n4074) );
  AN2 U1907 ( .A(n3645), .B(n4076), .Z(n3860) );
  OR2 U1908 ( .A(n4077), .B(n3727), .Z(n4076) );
  OR2 U1909 ( .A(n3918), .B(n3689), .Z(n4077) );
  OR2 U1910 ( .A(n3732), .B(n4078), .Z(n3689) );
  OR2 U1911 ( .A(n3947), .B(n3646), .Z(n4078) );
  IV U1912 ( .A(n1455), .Z(n3645) );
  AN2 U1913 ( .A(n4079), .B(n3954), .Z(n4069) );
  IV U1914 ( .A(n1449), .Z(n3954) );
  OR2 U1915 ( .A(n4080), .B(n4081), .Z(n4000) );
  OR2 U1916 ( .A(n4082), .B(n4083), .Z(n4081) );
  AN2 U1917 ( .A(U47_DATA121_0), .B(n4084), .Z(n4083) );
  OR2 U1918 ( .A(n4085), .B(n4024), .Z(n4084) );
  AN2 U1919 ( .A(n4086), .B(n3531), .Z(n4082) );
  AN2 U1920 ( .A(n4087), .B(n4088), .Z(n4080) );
  OR2 U1921 ( .A(n3982), .B(n3972), .Z(n4087) );
  IV U1922 ( .A(n1348), .Z(n3972) );
  IV U1923 ( .A(n1381), .Z(n3982) );
  AN2 U1924 ( .A(n1919), .B(n2112), .Z(n3702) );
  OR2 U1925 ( .A(n4008), .B(n4089), .Z(U20_Z_0) );
  OR2 U1926 ( .A(n4090), .B(n4091), .Z(n4089) );
  AN2 U1927 ( .A(n4092), .B(n3528), .Z(n4091) );
  IV U1928 ( .A(n2112), .Z(n3528) );
  OR2 U1929 ( .A(n4093), .B(n4094), .Z(n4092) );
  OR2 U1930 ( .A(n4095), .B(n4096), .Z(n4094) );
  OR2 U1931 ( .A(n4019), .B(n4041), .Z(n4096) );
  OR2 U1932 ( .A(n4097), .B(n4098), .Z(n4041) );
  AN2 U1933 ( .A(n4099), .B(n3531), .Z(n4098) );
  OR2 U1934 ( .A(n4004), .B(n4032), .Z(n4099) );
  OR2 U1935 ( .A(n4100), .B(n4101), .Z(n4032) );
  AN2 U1936 ( .A(n4102), .B(n3984), .Z(n4101) );
  AN2 U1937 ( .A(n4103), .B(n3974), .Z(n4100) );
  OR2 U1938 ( .A(n4104), .B(n4105), .Z(n4004) );
  AN2 U1939 ( .A(n4106), .B(n3988), .Z(n4105) );
  AN2 U1940 ( .A(n4107), .B(n3968), .Z(n4104) );
  AN2 U1941 ( .A(U47_DATA121_0), .B(n4030), .Z(n4097) );
  OR2 U1942 ( .A(n4108), .B(n4109), .Z(n4030) );
  AN2 U1943 ( .A(n4106), .B(n3984), .Z(n4109) );
  IV U1944 ( .A(n1248), .Z(n3984) );
  AN2 U1945 ( .A(n4107), .B(n3974), .Z(n4108) );
  IV U1946 ( .A(n1214), .Z(n3974) );
  OR2 U1947 ( .A(n4110), .B(n4003), .Z(n4019) );
  AN2 U1948 ( .A(U47_DATA121_0), .B(n4045), .Z(n4003) );
  OR2 U1949 ( .A(n4111), .B(n4112), .Z(n4045) );
  AN2 U1950 ( .A(n4102), .B(n3985), .Z(n4112) );
  AN2 U1951 ( .A(n4103), .B(n3971), .Z(n4111) );
  AN2 U1952 ( .A(n4113), .B(n4088), .Z(n4110) );
  OR2 U1953 ( .A(n3986), .B(n3973), .Z(n4113) );
  IV U1954 ( .A(n1146), .Z(n3973) );
  IV U1955 ( .A(n1179), .Z(n3986) );
  OR2 U1956 ( .A(n4114), .B(n4115), .Z(n4095) );
  AN2 U1957 ( .A(n4116), .B(n3531), .Z(n4115) );
  IV U1958 ( .A(U47_DATA121_0), .Z(n3531) );
  OR2 U1959 ( .A(n4024), .B(n4031), .Z(n4116) );
  OR2 U1960 ( .A(n4117), .B(n4118), .Z(n4031) );
  AN2 U1961 ( .A(n4106), .B(n3985), .Z(n4118) );
  IV U1962 ( .A(n1315), .Z(n3985) );
  AN2 U1963 ( .A(n4107), .B(n3971), .Z(n4117) );
  IV U1964 ( .A(n1282), .Z(n3971) );
  OR2 U1965 ( .A(n4119), .B(n4120), .Z(n4107) );
  OR2 U1966 ( .A(n4121), .B(n4122), .Z(n4024) );
  OR2 U1967 ( .A(n4123), .B(n3929), .Z(n4122) );
  AN2 U1968 ( .A(n1579), .B(n1578), .Z(n3929) );
  AN2 U1969 ( .A(n4079), .B(n3915), .Z(n4123) );
  IV U1970 ( .A(n1485), .Z(n3915) );
  OR2 U1971 ( .A(n3882), .B(n3916), .Z(n4079) );
  OR2 U1972 ( .A(n4124), .B(n4125), .Z(n4121) );
  AN2 U1973 ( .A(n4126), .B(n3887), .Z(n4125) );
  OR2 U1974 ( .A(n4127), .B(n4128), .Z(n4126) );
  OR2 U1975 ( .A(n3888), .B(n3881), .Z(n4128) );
  IV U1976 ( .A(n1536), .Z(n3881) );
  OR2 U1977 ( .A(n3947), .B(n3918), .Z(n4127) );
  IV U1978 ( .A(n1503), .Z(n3918) );
  IV U1979 ( .A(n1496), .Z(n3947) );
  AN2 U1980 ( .A(n4129), .B(n3951), .Z(n4124) );
  OR2 U1981 ( .A(n3882), .B(n4075), .Z(n4129) );
  OR2 U1982 ( .A(n3888), .B(n4130), .Z(n4075) );
  OR2 U1983 ( .A(n4059), .B(n3900), .Z(n4130) );
  OR2 U1984 ( .A(n3787), .B(n4131), .Z(n4059) );
  OR2 U1985 ( .A(n3791), .B(n3795), .Z(n4131) );
  IV U1986 ( .A(n1568), .Z(n3795) );
  IV U1987 ( .A(n1563), .Z(n3791) );
  IV U1988 ( .A(n1571), .Z(n3787) );
  IV U1989 ( .A(n1517), .Z(n3888) );
  AN2 U1990 ( .A(U47_DATA121_0), .B(n4025), .Z(n4114) );
  OR2 U1991 ( .A(n4085), .B(n4086), .Z(n4025) );
  OR2 U1992 ( .A(n4132), .B(n4133), .Z(n4086) );
  OR2 U1993 ( .A(n3847), .B(n4134), .Z(n4133) );
  OR2 U1994 ( .A(n3443), .B(n4135), .Z(n4134) );
  AN2 U1995 ( .A(n4136), .B(n3887), .Z(n4135) );
  IV U1996 ( .A(n1495), .Z(n3887) );
  OR2 U1997 ( .A(n4137), .B(n4138), .Z(n4136) );
  OR2 U1998 ( .A(n3900), .B(n4073), .Z(n4138) );
  OR2 U1999 ( .A(n3829), .B(n4139), .Z(n4073) );
  OR2 U2000 ( .A(n3851), .B(n3855), .Z(n4139) );
  IV U2001 ( .A(n1513), .Z(n3900) );
  OR2 U2002 ( .A(n3727), .B(n4140), .Z(n4137) );
  OR2 U2003 ( .A(n3646), .B(n3732), .Z(n4140) );
  AN2 U2004 ( .A(n3951), .B(n3829), .Z(n3443) );
  IV U2005 ( .A(n1528), .Z(n3829) );
  AN2 U2006 ( .A(n3646), .B(n3951), .Z(n3847) );
  IV U2007 ( .A(n1499), .Z(n3646) );
  OR2 U2008 ( .A(n4141), .B(n4142), .Z(n4132) );
  OR2 U2009 ( .A(n3447), .B(n3446), .Z(n4142) );
  AN2 U2010 ( .A(n3951), .B(n3855), .Z(n3446) );
  IV U2011 ( .A(n1523), .Z(n3855) );
  AN2 U2012 ( .A(n3951), .B(n3732), .Z(n3447) );
  IV U2013 ( .A(n1509), .Z(n3732) );
  OR2 U2014 ( .A(n3451), .B(n3450), .Z(n4141) );
  AN2 U2015 ( .A(n3951), .B(n3851), .Z(n3450) );
  IV U2016 ( .A(n1520), .Z(n3851) );
  AN2 U2017 ( .A(n3951), .B(n3727), .Z(n3451) );
  IV U2018 ( .A(n1506), .Z(n3727) );
  OR2 U2019 ( .A(n3937), .B(n4143), .Z(n4085) );
  OR2 U2020 ( .A(n4144), .B(n4145), .Z(n4143) );
  AN2 U2021 ( .A(n4102), .B(n3988), .Z(n4145) );
  IV U2022 ( .A(n1043), .Z(n3988) );
  AN2 U2023 ( .A(n4146), .B(n3968), .Z(n4144) );
  IV U2024 ( .A(n993), .Z(n3968) );
  OR2 U2025 ( .A(n4147), .B(n4061), .Z(n4146) );
  AN2 U2026 ( .A(n988), .B(n987), .Z(n3937) );
  OR2 U2027 ( .A(n4001), .B(n4148), .Z(n4093) );
  OR2 U2028 ( .A(n1643), .B(n4067), .Z(n4148) );
  AN2 U2029 ( .A(n3916), .B(n3951), .Z(n4067) );
  IV U2030 ( .A(n1540), .Z(n3951) );
  IV U2031 ( .A(n1489), .Z(n3916) );
  OR2 U2032 ( .A(n4149), .B(n4150), .Z(n4001) );
  OR2 U2033 ( .A(n3800), .B(n4151), .Z(n4150) );
  AN2 U2034 ( .A(n4152), .B(n3651), .Z(n4151) );
  OR2 U2035 ( .A(n3899), .B(n4153), .Z(n4152) );
  OR2 U2036 ( .A(n4103), .B(n4154), .Z(n4153) );
  OR2 U2037 ( .A(n4155), .B(n4061), .Z(n4103) );
  AN2 U2038 ( .A(n3651), .B(n4156), .Z(n3800) );
  OR2 U2039 ( .A(n4157), .B(n3725), .Z(n4156) );
  OR2 U2040 ( .A(n3831), .B(n3688), .Z(n4157) );
  OR2 U2041 ( .A(n3731), .B(n4158), .Z(n3688) );
  OR2 U2042 ( .A(n3856), .B(n3650), .Z(n4158) );
  IV U2043 ( .A(n1080), .Z(n3651) );
  AN2 U2044 ( .A(n4088), .B(n3989), .Z(n4149) );
  IV U2045 ( .A(n1113), .Z(n3989) );
  OR2 U2046 ( .A(n4102), .B(n4106), .Z(n4088) );
  OR2 U2047 ( .A(n4061), .B(n4119), .Z(n4106) );
  OR2 U2048 ( .A(n4154), .B(n4159), .Z(n4119) );
  OR2 U2049 ( .A(n3856), .B(n3831), .Z(n4159) );
  IV U2050 ( .A(n1031), .Z(n3831) );
  IV U2051 ( .A(n1026), .Z(n3856) );
  OR2 U2052 ( .A(n4160), .B(n4161), .Z(n4154) );
  OR2 U2053 ( .A(n3832), .B(n3852), .Z(n4161) );
  IV U2054 ( .A(n1023), .Z(n3852) );
  IV U2055 ( .A(n1012), .Z(n3832) );
  OR2 U2056 ( .A(n3848), .B(n3841), .Z(n4160) );
  IV U2057 ( .A(n1009), .Z(n3841) );
  IV U2058 ( .A(n1001), .Z(n3848) );
  OR2 U2059 ( .A(n3948), .B(n4162), .Z(n4061) );
  OR2 U2060 ( .A(n3944), .B(n3917), .Z(n4162) );
  IV U2061 ( .A(n994), .Z(n3917) );
  IV U2062 ( .A(n1006), .Z(n3944) );
  IV U2063 ( .A(n998), .Z(n3948) );
  OR2 U2064 ( .A(n4155), .B(n4120), .Z(n4102) );
  OR2 U2065 ( .A(n4163), .B(n4164), .Z(n4120) );
  OR2 U2066 ( .A(n3725), .B(n3899), .Z(n4164) );
  IV U2067 ( .A(n1016), .Z(n3899) );
  IV U2068 ( .A(n1072), .Z(n3725) );
  OR2 U2069 ( .A(n3650), .B(n3731), .Z(n4163) );
  IV U2070 ( .A(n1075), .Z(n3731) );
  IV U2071 ( .A(n1067), .Z(n3650) );
  OR2 U2072 ( .A(n4147), .B(n3882), .Z(n4155) );
  IV U2073 ( .A(n1044), .Z(n3882) );
  OR2 U2074 ( .A(n3890), .B(n3880), .Z(n4147) );
  IV U2075 ( .A(n1039), .Z(n3880) );
  IV U2076 ( .A(n1020), .Z(n3890) );
  AN2 U2077 ( .A(n1916), .B(n2112), .Z(n4090) );
  AN2 U2078 ( .A(n3594), .B(n3994), .Z(n4008) );
  OR2 U2079 ( .A(n3743), .B(n4036), .Z(n3994) );
  OR2 U2080 ( .A(n3660), .B(n3693), .Z(n4036) );
  OR2 U2081 ( .A(n3662), .B(n3657), .Z(n3693) );
  AN2 U2082 ( .A(n4165), .B(n3738), .Z(n3657) );
  IV U2083 ( .A(n1607), .Z(n4165) );
  AN2 U2084 ( .A(n4015), .B(n4014), .Z(n3662) );
  IV U2085 ( .A(n1594), .Z(n4014) );
  IV U2086 ( .A(n1601), .Z(n4015) );
  AN2 U2087 ( .A(n4166), .B(n3738), .Z(n3660) );
  IV U2088 ( .A(n1606), .Z(n3738) );
  OR2 U2089 ( .A(n3744), .B(n3739), .Z(n4166) );
  IV U2090 ( .A(n1616), .Z(n3739) );
  IV U2091 ( .A(n1610), .Z(n3744) );
  AN2 U2092 ( .A(n1591), .B(n1590), .Z(n3743) );
  AN2 U2093 ( .A(U47_DATA121_0), .B(n2112), .Z(n3594) );
endmodule

